// This is the unpowered netlist.
module wb_lfsr (i_clk,
    i_reset,
    i_wb_cyc,
    i_wb_stb,
    i_wb_we,
    o_wb_ack,
    o_wb_data,
    o_wb_stall,
    i_wb_addr,
    i_wb_data);
 input i_clk;
 input i_reset;
 input i_wb_cyc;
 input i_wb_stb;
 input i_wb_we;
 output o_wb_ack;
 output o_wb_data;
 output o_wb_stall;
 input [2:0] i_wb_addr;
 input [7:0] i_wb_data;

 wire net28;
 wire \FLSR_instance.flip_flop_instance[0].in ;
 wire \FLSR_instance.flip_flop_instance[0].out ;
 wire \FLSR_instance.flip_flop_instance[0].reset ;
 wire \FLSR_instance.flip_flop_instance[10].in ;
 wire \FLSR_instance.flip_flop_instance[10].out ;
 wire \FLSR_instance.flip_flop_instance[11].in ;
 wire \FLSR_instance.flip_flop_instance[11].out ;
 wire \FLSR_instance.flip_flop_instance[12].in ;
 wire \FLSR_instance.flip_flop_instance[12].out ;
 wire \FLSR_instance.flip_flop_instance[13].in ;
 wire \FLSR_instance.flip_flop_instance[13].out ;
 wire \FLSR_instance.flip_flop_instance[14].in ;
 wire \FLSR_instance.flip_flop_instance[14].out ;
 wire \FLSR_instance.flip_flop_instance[15].in ;
 wire \FLSR_instance.flip_flop_instance[15].out ;
 wire \FLSR_instance.flip_flop_instance[16].in ;
 wire \FLSR_instance.flip_flop_instance[16].out ;
 wire \FLSR_instance.flip_flop_instance[17].in ;
 wire \FLSR_instance.flip_flop_instance[17].out ;
 wire \FLSR_instance.flip_flop_instance[18].in ;
 wire \FLSR_instance.flip_flop_instance[18].out ;
 wire \FLSR_instance.flip_flop_instance[19].in ;
 wire \FLSR_instance.flip_flop_instance[19].out ;
 wire \FLSR_instance.flip_flop_instance[1].in ;
 wire \FLSR_instance.flip_flop_instance[1].out ;
 wire \FLSR_instance.flip_flop_instance[20].in ;
 wire \FLSR_instance.flip_flop_instance[20].out ;
 wire \FLSR_instance.flip_flop_instance[21].in ;
 wire \FLSR_instance.flip_flop_instance[21].out ;
 wire \FLSR_instance.flip_flop_instance[22].in ;
 wire \FLSR_instance.flip_flop_instance[22].out ;
 wire \FLSR_instance.flip_flop_instance[23].in ;
 wire \FLSR_instance.flip_flop_instance[23].out ;
 wire \FLSR_instance.flip_flop_instance[24].in ;
 wire \FLSR_instance.flip_flop_instance[24].out ;
 wire \FLSR_instance.flip_flop_instance[25].in ;
 wire \FLSR_instance.flip_flop_instance[25].out ;
 wire \FLSR_instance.flip_flop_instance[26].in ;
 wire \FLSR_instance.flip_flop_instance[26].out ;
 wire \FLSR_instance.flip_flop_instance[27].in ;
 wire \FLSR_instance.flip_flop_instance[27].out ;
 wire \FLSR_instance.flip_flop_instance[28].in ;
 wire \FLSR_instance.flip_flop_instance[28].out ;
 wire \FLSR_instance.flip_flop_instance[29].in ;
 wire \FLSR_instance.flip_flop_instance[29].out ;
 wire \FLSR_instance.flip_flop_instance[2].in ;
 wire \FLSR_instance.flip_flop_instance[2].out ;
 wire \FLSR_instance.flip_flop_instance[30].in ;
 wire \FLSR_instance.flip_flop_instance[30].out ;
 wire \FLSR_instance.flip_flop_instance[31].in ;
 wire \FLSR_instance.flip_flop_instance[31].out ;
 wire \FLSR_instance.flip_flop_instance[3].in ;
 wire \FLSR_instance.flip_flop_instance[3].out ;
 wire \FLSR_instance.flip_flop_instance[4].in ;
 wire \FLSR_instance.flip_flop_instance[4].out ;
 wire \FLSR_instance.flip_flop_instance[5].in ;
 wire \FLSR_instance.flip_flop_instance[5].out ;
 wire \FLSR_instance.flip_flop_instance[6].in ;
 wire \FLSR_instance.flip_flop_instance[6].out ;
 wire \FLSR_instance.flip_flop_instance[7].in ;
 wire \FLSR_instance.flip_flop_instance[7].out ;
 wire \FLSR_instance.flip_flop_instance[8].in ;
 wire \FLSR_instance.flip_flop_instance[8].out ;
 wire \FLSR_instance.flip_flop_instance[9].in ;
 wire \FLSR_instance.flip_flop_instance[9].out ;
 wire \FLSR_instance.load_seed ;
 wire \FLSR_instance.muxes[0].input_a ;
 wire \FLSR_instance.muxes[10].input_a ;
 wire \FLSR_instance.muxes[11].input_a ;
 wire \FLSR_instance.muxes[12].input_a ;
 wire \FLSR_instance.muxes[13].input_a ;
 wire \FLSR_instance.muxes[14].input_a ;
 wire \FLSR_instance.muxes[15].input_a ;
 wire \FLSR_instance.muxes[16].input_a ;
 wire \FLSR_instance.muxes[17].input_a ;
 wire \FLSR_instance.muxes[18].input_a ;
 wire \FLSR_instance.muxes[19].input_a ;
 wire \FLSR_instance.muxes[1].input_a ;
 wire \FLSR_instance.muxes[20].input_a ;
 wire \FLSR_instance.muxes[21].input_a ;
 wire \FLSR_instance.muxes[22].input_a ;
 wire \FLSR_instance.muxes[23].input_a ;
 wire \FLSR_instance.muxes[24].input_a ;
 wire \FLSR_instance.muxes[25].input_a ;
 wire \FLSR_instance.muxes[26].input_a ;
 wire \FLSR_instance.muxes[27].input_a ;
 wire \FLSR_instance.muxes[28].input_a ;
 wire \FLSR_instance.muxes[29].input_a ;
 wire \FLSR_instance.muxes[2].input_a ;
 wire \FLSR_instance.muxes[30].input_a ;
 wire \FLSR_instance.muxes[31].input_a ;
 wire \FLSR_instance.muxes[3].input_a ;
 wire \FLSR_instance.muxes[4].input_a ;
 wire \FLSR_instance.muxes[5].input_a ;
 wire \FLSR_instance.muxes[6].input_a ;
 wire \FLSR_instance.muxes[7].input_a ;
 wire \FLSR_instance.muxes[8].input_a ;
 wire \FLSR_instance.muxes[9].input_a ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net11));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_82 ();
 sky130_fd_sc_hd__clkbuf_4 _167_ (.A(\FLSR_instance.load_seed ),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _168_ (.A0(\FLSR_instance.flip_flop_instance[30].out ),
    .A1(\FLSR_instance.muxes[31].input_a ),
    .S(_068_),
    .X(_069_));
 sky130_fd_sc_hd__clkbuf_1 _169_ (.A(_069_),
    .X(\FLSR_instance.flip_flop_instance[31].in ));
 sky130_fd_sc_hd__mux2_1 _170_ (.A0(\FLSR_instance.flip_flop_instance[29].out ),
    .A1(\FLSR_instance.muxes[30].input_a ),
    .S(_068_),
    .X(_070_));
 sky130_fd_sc_hd__clkbuf_1 _171_ (.A(_070_),
    .X(\FLSR_instance.flip_flop_instance[30].in ));
 sky130_fd_sc_hd__mux2_1 _172_ (.A0(\FLSR_instance.flip_flop_instance[28].out ),
    .A1(\FLSR_instance.muxes[29].input_a ),
    .S(_068_),
    .X(_071_));
 sky130_fd_sc_hd__clkbuf_1 _173_ (.A(_071_),
    .X(\FLSR_instance.flip_flop_instance[29].in ));
 sky130_fd_sc_hd__mux2_1 _174_ (.A0(\FLSR_instance.flip_flop_instance[27].out ),
    .A1(\FLSR_instance.muxes[28].input_a ),
    .S(_068_),
    .X(_072_));
 sky130_fd_sc_hd__clkbuf_1 _175_ (.A(_072_),
    .X(\FLSR_instance.flip_flop_instance[28].in ));
 sky130_fd_sc_hd__mux2_1 _176_ (.A0(\FLSR_instance.flip_flop_instance[26].out ),
    .A1(\FLSR_instance.muxes[27].input_a ),
    .S(_068_),
    .X(_073_));
 sky130_fd_sc_hd__clkbuf_1 _177_ (.A(_073_),
    .X(\FLSR_instance.flip_flop_instance[27].in ));
 sky130_fd_sc_hd__mux2_1 _178_ (.A0(\FLSR_instance.flip_flop_instance[25].out ),
    .A1(\FLSR_instance.muxes[26].input_a ),
    .S(_068_),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _179_ (.A(_074_),
    .X(\FLSR_instance.flip_flop_instance[26].in ));
 sky130_fd_sc_hd__mux2_1 _180_ (.A0(\FLSR_instance.flip_flop_instance[24].out ),
    .A1(\FLSR_instance.muxes[25].input_a ),
    .S(_068_),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _181_ (.A(_075_),
    .X(\FLSR_instance.flip_flop_instance[25].in ));
 sky130_fd_sc_hd__mux2_1 _182_ (.A0(\FLSR_instance.flip_flop_instance[23].out ),
    .A1(\FLSR_instance.muxes[24].input_a ),
    .S(_068_),
    .X(_076_));
 sky130_fd_sc_hd__clkbuf_1 _183_ (.A(_076_),
    .X(\FLSR_instance.flip_flop_instance[24].in ));
 sky130_fd_sc_hd__mux2_1 _184_ (.A0(\FLSR_instance.flip_flop_instance[22].out ),
    .A1(\FLSR_instance.muxes[23].input_a ),
    .S(_068_),
    .X(_077_));
 sky130_fd_sc_hd__clkbuf_1 _185_ (.A(_077_),
    .X(\FLSR_instance.flip_flop_instance[23].in ));
 sky130_fd_sc_hd__clkbuf_4 _186_ (.A(\FLSR_instance.load_seed ),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _187_ (.A0(\FLSR_instance.flip_flop_instance[21].out ),
    .A1(\FLSR_instance.muxes[22].input_a ),
    .S(_078_),
    .X(_079_));
 sky130_fd_sc_hd__clkbuf_1 _188_ (.A(_079_),
    .X(\FLSR_instance.flip_flop_instance[22].in ));
 sky130_fd_sc_hd__mux2_1 _189_ (.A0(\FLSR_instance.flip_flop_instance[20].out ),
    .A1(\FLSR_instance.muxes[21].input_a ),
    .S(_078_),
    .X(_080_));
 sky130_fd_sc_hd__clkbuf_1 _190_ (.A(_080_),
    .X(\FLSR_instance.flip_flop_instance[21].in ));
 sky130_fd_sc_hd__mux2_1 _191_ (.A0(\FLSR_instance.flip_flop_instance[19].out ),
    .A1(\FLSR_instance.muxes[20].input_a ),
    .S(_078_),
    .X(_081_));
 sky130_fd_sc_hd__clkbuf_1 _192_ (.A(_081_),
    .X(\FLSR_instance.flip_flop_instance[20].in ));
 sky130_fd_sc_hd__mux2_1 _193_ (.A0(\FLSR_instance.flip_flop_instance[18].out ),
    .A1(\FLSR_instance.muxes[19].input_a ),
    .S(_078_),
    .X(_082_));
 sky130_fd_sc_hd__clkbuf_1 _194_ (.A(_082_),
    .X(\FLSR_instance.flip_flop_instance[19].in ));
 sky130_fd_sc_hd__mux2_1 _195_ (.A0(\FLSR_instance.flip_flop_instance[17].out ),
    .A1(\FLSR_instance.muxes[18].input_a ),
    .S(_078_),
    .X(_083_));
 sky130_fd_sc_hd__clkbuf_1 _196_ (.A(_083_),
    .X(\FLSR_instance.flip_flop_instance[18].in ));
 sky130_fd_sc_hd__mux2_1 _197_ (.A0(\FLSR_instance.flip_flop_instance[16].out ),
    .A1(\FLSR_instance.muxes[17].input_a ),
    .S(_078_),
    .X(_084_));
 sky130_fd_sc_hd__clkbuf_1 _198_ (.A(_084_),
    .X(\FLSR_instance.flip_flop_instance[17].in ));
 sky130_fd_sc_hd__mux2_1 _199_ (.A0(\FLSR_instance.flip_flop_instance[15].out ),
    .A1(\FLSR_instance.muxes[16].input_a ),
    .S(_078_),
    .X(_085_));
 sky130_fd_sc_hd__clkbuf_1 _200_ (.A(_085_),
    .X(\FLSR_instance.flip_flop_instance[16].in ));
 sky130_fd_sc_hd__mux2_1 _201_ (.A0(\FLSR_instance.flip_flop_instance[14].out ),
    .A1(\FLSR_instance.muxes[15].input_a ),
    .S(_078_),
    .X(_086_));
 sky130_fd_sc_hd__clkbuf_1 _202_ (.A(_086_),
    .X(\FLSR_instance.flip_flop_instance[15].in ));
 sky130_fd_sc_hd__mux2_1 _203_ (.A0(\FLSR_instance.flip_flop_instance[13].out ),
    .A1(\FLSR_instance.muxes[14].input_a ),
    .S(_078_),
    .X(_087_));
 sky130_fd_sc_hd__clkbuf_1 _204_ (.A(_087_),
    .X(\FLSR_instance.flip_flop_instance[14].in ));
 sky130_fd_sc_hd__mux2_1 _205_ (.A0(\FLSR_instance.flip_flop_instance[12].out ),
    .A1(\FLSR_instance.muxes[13].input_a ),
    .S(_078_),
    .X(_088_));
 sky130_fd_sc_hd__clkbuf_1 _206_ (.A(_088_),
    .X(\FLSR_instance.flip_flop_instance[13].in ));
 sky130_fd_sc_hd__clkbuf_4 _207_ (.A(\FLSR_instance.load_seed ),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _208_ (.A0(\FLSR_instance.flip_flop_instance[11].out ),
    .A1(\FLSR_instance.muxes[12].input_a ),
    .S(_089_),
    .X(_090_));
 sky130_fd_sc_hd__clkbuf_1 _209_ (.A(_090_),
    .X(\FLSR_instance.flip_flop_instance[12].in ));
 sky130_fd_sc_hd__mux2_1 _210_ (.A0(\FLSR_instance.flip_flop_instance[10].out ),
    .A1(\FLSR_instance.muxes[11].input_a ),
    .S(_089_),
    .X(_091_));
 sky130_fd_sc_hd__clkbuf_1 _211_ (.A(_091_),
    .X(\FLSR_instance.flip_flop_instance[11].in ));
 sky130_fd_sc_hd__mux2_1 _212_ (.A0(\FLSR_instance.flip_flop_instance[9].out ),
    .A1(\FLSR_instance.muxes[10].input_a ),
    .S(_089_),
    .X(_092_));
 sky130_fd_sc_hd__clkbuf_1 _213_ (.A(_092_),
    .X(\FLSR_instance.flip_flop_instance[10].in ));
 sky130_fd_sc_hd__mux2_1 _214_ (.A0(\FLSR_instance.flip_flop_instance[8].out ),
    .A1(\FLSR_instance.muxes[9].input_a ),
    .S(_089_),
    .X(_093_));
 sky130_fd_sc_hd__clkbuf_1 _215_ (.A(_093_),
    .X(\FLSR_instance.flip_flop_instance[9].in ));
 sky130_fd_sc_hd__mux2_1 _216_ (.A0(\FLSR_instance.flip_flop_instance[7].out ),
    .A1(\FLSR_instance.muxes[8].input_a ),
    .S(_089_),
    .X(_094_));
 sky130_fd_sc_hd__clkbuf_1 _217_ (.A(_094_),
    .X(\FLSR_instance.flip_flop_instance[8].in ));
 sky130_fd_sc_hd__mux2_1 _218_ (.A0(\FLSR_instance.flip_flop_instance[6].out ),
    .A1(\FLSR_instance.muxes[7].input_a ),
    .S(_089_),
    .X(_095_));
 sky130_fd_sc_hd__clkbuf_1 _219_ (.A(_095_),
    .X(\FLSR_instance.flip_flop_instance[7].in ));
 sky130_fd_sc_hd__mux2_1 _220_ (.A0(\FLSR_instance.flip_flop_instance[5].out ),
    .A1(\FLSR_instance.muxes[6].input_a ),
    .S(_089_),
    .X(_096_));
 sky130_fd_sc_hd__clkbuf_1 _221_ (.A(_096_),
    .X(\FLSR_instance.flip_flop_instance[6].in ));
 sky130_fd_sc_hd__mux2_1 _222_ (.A0(\FLSR_instance.flip_flop_instance[4].out ),
    .A1(\FLSR_instance.muxes[5].input_a ),
    .S(_089_),
    .X(_097_));
 sky130_fd_sc_hd__clkbuf_1 _223_ (.A(_097_),
    .X(\FLSR_instance.flip_flop_instance[5].in ));
 sky130_fd_sc_hd__mux2_1 _224_ (.A0(\FLSR_instance.flip_flop_instance[3].out ),
    .A1(\FLSR_instance.muxes[4].input_a ),
    .S(_089_),
    .X(_098_));
 sky130_fd_sc_hd__clkbuf_1 _225_ (.A(_098_),
    .X(\FLSR_instance.flip_flop_instance[4].in ));
 sky130_fd_sc_hd__mux2_1 _226_ (.A0(\FLSR_instance.flip_flop_instance[2].out ),
    .A1(\FLSR_instance.muxes[3].input_a ),
    .S(_089_),
    .X(_099_));
 sky130_fd_sc_hd__clkbuf_1 _227_ (.A(_099_),
    .X(\FLSR_instance.flip_flop_instance[3].in ));
 sky130_fd_sc_hd__mux2_1 _228_ (.A0(\FLSR_instance.flip_flop_instance[1].out ),
    .A1(\FLSR_instance.muxes[2].input_a ),
    .S(\FLSR_instance.load_seed ),
    .X(_100_));
 sky130_fd_sc_hd__clkbuf_1 _229_ (.A(_100_),
    .X(\FLSR_instance.flip_flop_instance[2].in ));
 sky130_fd_sc_hd__mux2_1 _230_ (.A0(\FLSR_instance.flip_flop_instance[0].out ),
    .A1(\FLSR_instance.muxes[1].input_a ),
    .S(\FLSR_instance.load_seed ),
    .X(_101_));
 sky130_fd_sc_hd__clkbuf_1 _231_ (.A(_101_),
    .X(\FLSR_instance.flip_flop_instance[1].in ));
 sky130_fd_sc_hd__xor2_1 _232_ (.A(\FLSR_instance.flip_flop_instance[6].out ),
    .B(\FLSR_instance.flip_flop_instance[31].out ),
    .X(_102_));
 sky130_fd_sc_hd__xnor2_1 _233_ (.A(\FLSR_instance.flip_flop_instance[5].out ),
    .B(\FLSR_instance.flip_flop_instance[1].out ),
    .Y(_103_));
 sky130_fd_sc_hd__xnor2_1 _234_ (.A(_102_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__mux2_1 _235_ (.A0(_104_),
    .A1(\FLSR_instance.muxes[0].input_a ),
    .S(\FLSR_instance.load_seed ),
    .X(_105_));
 sky130_fd_sc_hd__clkbuf_1 _236_ (.A(_105_),
    .X(\FLSR_instance.flip_flop_instance[0].in ));
 sky130_fd_sc_hd__and3b_2 _237_ (.A_N(net5),
    .B(net4),
    .C(net3),
    .X(_106_));
 sky130_fd_sc_hd__and2_1 _238_ (.A(net7),
    .B(_106_),
    .X(_107_));
 sky130_fd_sc_hd__and3_1 _239_ (.A(net15),
    .B(net16),
    .C(net6),
    .X(_108_));
 sky130_fd_sc_hd__or3b_2 _240_ (.A(net4),
    .B(net3),
    .C_N(net5),
    .X(_109_));
 sky130_fd_sc_hd__or3b_1 _241_ (.A(net5),
    .B(net3),
    .C_N(net4),
    .X(_110_));
 sky130_fd_sc_hd__o2111a_4 _242_ (.A1(net5),
    .A2(net4),
    .B1(_108_),
    .C1(_109_),
    .D1(_110_),
    .X(_111_));
 sky130_fd_sc_hd__mux2_1 _243_ (.A0(\FLSR_instance.muxes[24].input_a ),
    .A1(_107_),
    .S(_111_),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_1 _244_ (.A(_112_),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _245_ (.A(net8),
    .B(_106_),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _246_ (.A0(\FLSR_instance.muxes[25].input_a ),
    .A1(_113_),
    .S(_111_),
    .X(_114_));
 sky130_fd_sc_hd__clkbuf_1 _247_ (.A(_114_),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _248_ (.A(net9),
    .B(_106_),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _249_ (.A0(\FLSR_instance.muxes[26].input_a ),
    .A1(_115_),
    .S(_111_),
    .X(_116_));
 sky130_fd_sc_hd__clkbuf_1 _250_ (.A(_116_),
    .X(_034_));
 sky130_fd_sc_hd__and2_1 _251_ (.A(net10),
    .B(_106_),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _252_ (.A0(\FLSR_instance.muxes[27].input_a ),
    .A1(_117_),
    .S(_111_),
    .X(_118_));
 sky130_fd_sc_hd__clkbuf_1 _253_ (.A(_118_),
    .X(_035_));
 sky130_fd_sc_hd__and2_1 _254_ (.A(net11),
    .B(_106_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _255_ (.A0(\FLSR_instance.muxes[28].input_a ),
    .A1(_119_),
    .S(_111_),
    .X(_120_));
 sky130_fd_sc_hd__clkbuf_1 _256_ (.A(_120_),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _257_ (.A(net12),
    .B(_106_),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _258_ (.A0(\FLSR_instance.muxes[29].input_a ),
    .A1(_121_),
    .S(_111_),
    .X(_122_));
 sky130_fd_sc_hd__clkbuf_1 _259_ (.A(_122_),
    .X(_037_));
 sky130_fd_sc_hd__and2_1 _260_ (.A(net13),
    .B(_106_),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _261_ (.A0(\FLSR_instance.muxes[30].input_a ),
    .A1(_123_),
    .S(_111_),
    .X(_124_));
 sky130_fd_sc_hd__clkbuf_1 _262_ (.A(_124_),
    .X(_038_));
 sky130_fd_sc_hd__and2_1 _263_ (.A(net14),
    .B(_106_),
    .X(_125_));
 sky130_fd_sc_hd__mux2_1 _264_ (.A0(\FLSR_instance.muxes[31].input_a ),
    .A1(_125_),
    .S(_111_),
    .X(_126_));
 sky130_fd_sc_hd__clkbuf_1 _265_ (.A(_126_),
    .X(_039_));
 sky130_fd_sc_hd__inv_2 _266_ (.A(net3),
    .Y(_127_));
 sky130_fd_sc_hd__o2111a_1 _267_ (.A1(net4),
    .A2(net3),
    .B1(net15),
    .C1(net16),
    .D1(net6),
    .X(_128_));
 sky130_fd_sc_hd__o21ai_4 _268_ (.A1(net5),
    .A2(_127_),
    .B1(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__and2b_1 _269_ (.A_N(net5),
    .B(net4),
    .X(_130_));
 sky130_fd_sc_hd__and3_1 _270_ (.A(_127_),
    .B(_130_),
    .C(_128_),
    .X(_131_));
 sky130_fd_sc_hd__buf_2 _271_ (.A(_131_),
    .X(_132_));
 sky130_fd_sc_hd__a22o_1 _272_ (.A1(\FLSR_instance.muxes[16].input_a ),
    .A2(_129_),
    .B1(_132_),
    .B2(net7),
    .X(_040_));
 sky130_fd_sc_hd__a22o_1 _273_ (.A1(\FLSR_instance.muxes[17].input_a ),
    .A2(_129_),
    .B1(_132_),
    .B2(net8),
    .X(_041_));
 sky130_fd_sc_hd__a22o_1 _274_ (.A1(\FLSR_instance.muxes[18].input_a ),
    .A2(_129_),
    .B1(_132_),
    .B2(net9),
    .X(_042_));
 sky130_fd_sc_hd__a22o_1 _275_ (.A1(\FLSR_instance.muxes[19].input_a ),
    .A2(_129_),
    .B1(_132_),
    .B2(net10),
    .X(_043_));
 sky130_fd_sc_hd__a22o_1 _276_ (.A1(\FLSR_instance.muxes[20].input_a ),
    .A2(_129_),
    .B1(_132_),
    .B2(net11),
    .X(_044_));
 sky130_fd_sc_hd__a22o_1 _277_ (.A1(\FLSR_instance.muxes[21].input_a ),
    .A2(_129_),
    .B1(_132_),
    .B2(net12),
    .X(_045_));
 sky130_fd_sc_hd__a22o_1 _278_ (.A1(\FLSR_instance.muxes[22].input_a ),
    .A2(_129_),
    .B1(_132_),
    .B2(net13),
    .X(_046_));
 sky130_fd_sc_hd__a22o_1 _279_ (.A1(\FLSR_instance.muxes[23].input_a ),
    .A2(_129_),
    .B1(_132_),
    .B2(net14),
    .X(_047_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(net8),
    .Y(_133_));
 sky130_fd_sc_hd__nor2_1 _281_ (.A(_133_),
    .B(_109_),
    .Y(_134_));
 sky130_fd_sc_hd__and2_1 _282_ (.A(net5),
    .B(_108_),
    .X(_135_));
 sky130_fd_sc_hd__mux2_1 _283_ (.A0(_068_),
    .A1(_134_),
    .S(_135_),
    .X(_136_));
 sky130_fd_sc_hd__clkbuf_1 _284_ (.A(_136_),
    .X(_048_));
 sky130_fd_sc_hd__nor3_2 _285_ (.A(net5),
    .B(net4),
    .C(net3),
    .Y(_137_));
 sky130_fd_sc_hd__and2_1 _286_ (.A(net7),
    .B(_137_),
    .X(_138_));
 sky130_fd_sc_hd__o2111a_4 _287_ (.A1(net5),
    .A2(_127_),
    .B1(_108_),
    .C1(_109_),
    .D1(_110_),
    .X(_139_));
 sky130_fd_sc_hd__mux2_1 _288_ (.A0(\FLSR_instance.muxes[0].input_a ),
    .A1(_138_),
    .S(_139_),
    .X(_140_));
 sky130_fd_sc_hd__clkbuf_1 _289_ (.A(_140_),
    .X(_049_));
 sky130_fd_sc_hd__and2_1 _290_ (.A(net8),
    .B(_137_),
    .X(_141_));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(\FLSR_instance.muxes[1].input_a ),
    .A1(_141_),
    .S(_139_),
    .X(_142_));
 sky130_fd_sc_hd__clkbuf_1 _292_ (.A(_142_),
    .X(_050_));
 sky130_fd_sc_hd__and2_1 _293_ (.A(net9),
    .B(_137_),
    .X(_143_));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(\FLSR_instance.muxes[2].input_a ),
    .A1(_143_),
    .S(_139_),
    .X(_144_));
 sky130_fd_sc_hd__clkbuf_1 _295_ (.A(_144_),
    .X(_051_));
 sky130_fd_sc_hd__and2_1 _296_ (.A(net10),
    .B(_137_),
    .X(_145_));
 sky130_fd_sc_hd__mux2_1 _297_ (.A0(\FLSR_instance.muxes[3].input_a ),
    .A1(_145_),
    .S(_139_),
    .X(_146_));
 sky130_fd_sc_hd__clkbuf_1 _298_ (.A(_146_),
    .X(_052_));
 sky130_fd_sc_hd__and2_1 _299_ (.A(net11),
    .B(_137_),
    .X(_147_));
 sky130_fd_sc_hd__mux2_1 _300_ (.A0(\FLSR_instance.muxes[4].input_a ),
    .A1(_147_),
    .S(_139_),
    .X(_148_));
 sky130_fd_sc_hd__clkbuf_1 _301_ (.A(_148_),
    .X(_053_));
 sky130_fd_sc_hd__and2_1 _302_ (.A(net12),
    .B(_137_),
    .X(_149_));
 sky130_fd_sc_hd__mux2_1 _303_ (.A0(\FLSR_instance.muxes[5].input_a ),
    .A1(_149_),
    .S(_139_),
    .X(_150_));
 sky130_fd_sc_hd__clkbuf_1 _304_ (.A(_150_),
    .X(_054_));
 sky130_fd_sc_hd__and2_1 _305_ (.A(net13),
    .B(_137_),
    .X(_151_));
 sky130_fd_sc_hd__mux2_1 _306_ (.A0(\FLSR_instance.muxes[6].input_a ),
    .A1(_151_),
    .S(_139_),
    .X(_152_));
 sky130_fd_sc_hd__clkbuf_1 _307_ (.A(_152_),
    .X(_055_));
 sky130_fd_sc_hd__and2_1 _308_ (.A(net14),
    .B(_137_),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _309_ (.A0(\FLSR_instance.muxes[7].input_a ),
    .A1(_153_),
    .S(_139_),
    .X(_154_));
 sky130_fd_sc_hd__clkbuf_1 _310_ (.A(_154_),
    .X(_056_));
 sky130_fd_sc_hd__or2b_1 _311_ (.A(_130_),
    .B_N(_128_),
    .X(_155_));
 sky130_fd_sc_hd__buf_2 _312_ (.A(_155_),
    .X(_156_));
 sky130_fd_sc_hd__and4bb_1 _313_ (.A_N(net5),
    .B_N(net4),
    .C(net3),
    .D(_128_),
    .X(_157_));
 sky130_fd_sc_hd__buf_2 _314_ (.A(_157_),
    .X(_158_));
 sky130_fd_sc_hd__a22o_1 _315_ (.A1(\FLSR_instance.muxes[8].input_a ),
    .A2(_156_),
    .B1(_158_),
    .B2(net7),
    .X(_057_));
 sky130_fd_sc_hd__a22o_1 _316_ (.A1(\FLSR_instance.muxes[9].input_a ),
    .A2(_156_),
    .B1(_158_),
    .B2(net8),
    .X(_058_));
 sky130_fd_sc_hd__a22o_1 _317_ (.A1(\FLSR_instance.muxes[10].input_a ),
    .A2(_156_),
    .B1(_158_),
    .B2(net9),
    .X(_059_));
 sky130_fd_sc_hd__a22o_1 _318_ (.A1(\FLSR_instance.muxes[11].input_a ),
    .A2(_156_),
    .B1(_158_),
    .B2(net10),
    .X(_060_));
 sky130_fd_sc_hd__a22o_1 _319_ (.A1(\FLSR_instance.muxes[12].input_a ),
    .A2(_156_),
    .B1(_158_),
    .B2(net11),
    .X(_061_));
 sky130_fd_sc_hd__a22o_1 _320_ (.A1(\FLSR_instance.muxes[13].input_a ),
    .A2(_156_),
    .B1(_158_),
    .B2(net12),
    .X(_062_));
 sky130_fd_sc_hd__a22o_1 _321_ (.A1(\FLSR_instance.muxes[14].input_a ),
    .A2(_156_),
    .B1(_158_),
    .B2(net13),
    .X(_063_));
 sky130_fd_sc_hd__a22o_1 _322_ (.A1(\FLSR_instance.muxes[15].input_a ),
    .A2(_156_),
    .B1(_158_),
    .B2(net14),
    .X(_064_));
 sky130_fd_sc_hd__and2b_1 _323_ (.A_N(net2),
    .B(net15),
    .X(_159_));
 sky130_fd_sc_hd__clkbuf_1 _324_ (.A(_159_),
    .X(_065_));
 sky130_fd_sc_hd__and3b_1 _325_ (.A_N(net16),
    .B(net6),
    .C(net15),
    .X(_160_));
 sky130_fd_sc_hd__mux2_1 _326_ (.A0(net18),
    .A1(_104_),
    .S(_160_),
    .X(_161_));
 sky130_fd_sc_hd__clkbuf_1 _327_ (.A(_161_),
    .X(_066_));
 sky130_fd_sc_hd__or3_1 _328_ (.A(net7),
    .B(net4),
    .C(net3),
    .X(_162_));
 sky130_fd_sc_hd__mux2_1 _329_ (.A0(\FLSR_instance.flip_flop_instance[0].reset ),
    .A1(_162_),
    .S(_135_),
    .X(_163_));
 sky130_fd_sc_hd__clkbuf_1 _330_ (.A(_163_),
    .X(_067_));
 sky130_fd_sc_hd__buf_4 _331_ (.A(\FLSR_instance.flip_flop_instance[0].reset ),
    .X(_164_));
 sky130_fd_sc_hd__inv_2 _332_ (.A(_164_),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _333_ (.A(_164_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _334_ (.A(_164_),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _335_ (.A(_164_),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _336_ (.A(_164_),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _337_ (.A(_164_),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _338_ (.A(_164_),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _339_ (.A(_164_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _340_ (.A(_164_),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _341_ (.A(_164_),
    .Y(_009_));
 sky130_fd_sc_hd__buf_4 _342_ (.A(\FLSR_instance.flip_flop_instance[0].reset ),
    .X(_165_));
 sky130_fd_sc_hd__inv_2 _343_ (.A(_165_),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _344_ (.A(_165_),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _345_ (.A(_165_),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _346_ (.A(_165_),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _347_ (.A(_165_),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _348_ (.A(_165_),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _349_ (.A(_165_),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _350_ (.A(_165_),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _351_ (.A(_165_),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _352_ (.A(_165_),
    .Y(_019_));
 sky130_fd_sc_hd__buf_4 _353_ (.A(\FLSR_instance.flip_flop_instance[0].reset ),
    .X(_166_));
 sky130_fd_sc_hd__inv_2 _354_ (.A(_166_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _355_ (.A(_166_),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _356_ (.A(_166_),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _357_ (.A(_166_),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _358_ (.A(_166_),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _359_ (.A(_166_),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _360_ (.A(_166_),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _361_ (.A(_166_),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _362_ (.A(_166_),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _363_ (.A(_166_),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _364_ (.A(\FLSR_instance.flip_flop_instance[0].reset ),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _365_ (.A(\FLSR_instance.flip_flop_instance[0].reset ),
    .Y(_031_));
 sky130_fd_sc_hd__dfxtp_1 _366_ (.CLK(net19),
    .D(_032_),
    .Q(\FLSR_instance.muxes[24].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _367_ (.CLK(net19),
    .D(_033_),
    .Q(\FLSR_instance.muxes[25].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _368_ (.CLK(net19),
    .D(_034_),
    .Q(\FLSR_instance.muxes[26].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _369_ (.CLK(net19),
    .D(_035_),
    .Q(\FLSR_instance.muxes[27].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _370_ (.CLK(net19),
    .D(_036_),
    .Q(\FLSR_instance.muxes[28].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _371_ (.CLK(net20),
    .D(_037_),
    .Q(\FLSR_instance.muxes[29].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _372_ (.CLK(net20),
    .D(_038_),
    .Q(\FLSR_instance.muxes[30].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _373_ (.CLK(net20),
    .D(_039_),
    .Q(\FLSR_instance.muxes[31].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _374_ (.CLK(net21),
    .D(_040_),
    .Q(\FLSR_instance.muxes[16].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _375_ (.CLK(net22),
    .D(_041_),
    .Q(\FLSR_instance.muxes[17].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _376_ (.CLK(net21),
    .D(_042_),
    .Q(\FLSR_instance.muxes[18].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _377_ (.CLK(net21),
    .D(_043_),
    .Q(\FLSR_instance.muxes[19].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _378_ (.CLK(net21),
    .D(_044_),
    .Q(\FLSR_instance.muxes[20].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _379_ (.CLK(net22),
    .D(_045_),
    .Q(\FLSR_instance.muxes[21].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _380_ (.CLK(net21),
    .D(_046_),
    .Q(\FLSR_instance.muxes[22].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _381_ (.CLK(net22),
    .D(_047_),
    .Q(\FLSR_instance.muxes[23].input_a ));
 sky130_fd_sc_hd__dfxtp_2 _382_ (.CLK(net23),
    .D(_048_),
    .Q(\FLSR_instance.load_seed ));
 sky130_fd_sc_hd__dfxtp_1 _383_ (.CLK(net23),
    .D(_049_),
    .Q(\FLSR_instance.muxes[0].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _384_ (.CLK(net23),
    .D(_050_),
    .Q(\FLSR_instance.muxes[1].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _385_ (.CLK(net24),
    .D(_051_),
    .Q(\FLSR_instance.muxes[2].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _386_ (.CLK(net24),
    .D(_052_),
    .Q(\FLSR_instance.muxes[3].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _387_ (.CLK(net25),
    .D(_053_),
    .Q(\FLSR_instance.muxes[4].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _388_ (.CLK(net24),
    .D(_054_),
    .Q(\FLSR_instance.muxes[5].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _389_ (.CLK(net23),
    .D(_055_),
    .Q(\FLSR_instance.muxes[6].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _390_ (.CLK(net23),
    .D(_056_),
    .Q(\FLSR_instance.muxes[7].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _391_ (.CLK(net25),
    .D(_057_),
    .Q(\FLSR_instance.muxes[8].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _392_ (.CLK(net25),
    .D(_058_),
    .Q(\FLSR_instance.muxes[9].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _393_ (.CLK(net25),
    .D(_059_),
    .Q(\FLSR_instance.muxes[10].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _394_ (.CLK(net26),
    .D(_060_),
    .Q(\FLSR_instance.muxes[11].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _395_ (.CLK(net25),
    .D(_061_),
    .Q(\FLSR_instance.muxes[12].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _396_ (.CLK(net25),
    .D(_062_),
    .Q(\FLSR_instance.muxes[13].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _397_ (.CLK(net25),
    .D(_063_),
    .Q(\FLSR_instance.muxes[14].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _398_ (.CLK(net22),
    .D(_064_),
    .Q(\FLSR_instance.muxes[15].input_a ));
 sky130_fd_sc_hd__dfxtp_1 _399_ (.CLK(net23),
    .D(_065_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _400_ (.CLK(net24),
    .D(_066_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_2 _401_ (.CLK(net25),
    .D(_067_),
    .Q(\FLSR_instance.flip_flop_instance[0].reset ));
 sky130_fd_sc_hd__dfrtp_1 _402_ (.CLK(net23),
    .D(\FLSR_instance.flip_flop_instance[31].in ),
    .RESET_B(_000_),
    .Q(\FLSR_instance.flip_flop_instance[31].out ));
 sky130_fd_sc_hd__dfrtp_1 _403_ (.CLK(net20),
    .D(\FLSR_instance.flip_flop_instance[30].in ),
    .RESET_B(_001_),
    .Q(\FLSR_instance.flip_flop_instance[30].out ));
 sky130_fd_sc_hd__dfrtp_1 _404_ (.CLK(net20),
    .D(\FLSR_instance.flip_flop_instance[29].in ),
    .RESET_B(_002_),
    .Q(\FLSR_instance.flip_flop_instance[29].out ));
 sky130_fd_sc_hd__dfrtp_1 _405_ (.CLK(net20),
    .D(\FLSR_instance.flip_flop_instance[28].in ),
    .RESET_B(_003_),
    .Q(\FLSR_instance.flip_flop_instance[28].out ));
 sky130_fd_sc_hd__dfrtp_1 _406_ (.CLK(net19),
    .D(\FLSR_instance.flip_flop_instance[27].in ),
    .RESET_B(_004_),
    .Q(\FLSR_instance.flip_flop_instance[27].out ));
 sky130_fd_sc_hd__dfrtp_1 _407_ (.CLK(net19),
    .D(\FLSR_instance.flip_flop_instance[26].in ),
    .RESET_B(_005_),
    .Q(\FLSR_instance.flip_flop_instance[26].out ));
 sky130_fd_sc_hd__dfrtp_1 _408_ (.CLK(net19),
    .D(\FLSR_instance.flip_flop_instance[25].in ),
    .RESET_B(_006_),
    .Q(\FLSR_instance.flip_flop_instance[25].out ));
 sky130_fd_sc_hd__dfrtp_1 _409_ (.CLK(net19),
    .D(\FLSR_instance.flip_flop_instance[24].in ),
    .RESET_B(_007_),
    .Q(\FLSR_instance.flip_flop_instance[24].out ));
 sky130_fd_sc_hd__dfrtp_1 _410_ (.CLK(net20),
    .D(\FLSR_instance.flip_flop_instance[23].in ),
    .RESET_B(_008_),
    .Q(\FLSR_instance.flip_flop_instance[23].out ));
 sky130_fd_sc_hd__dfrtp_1 _411_ (.CLK(net19),
    .D(\FLSR_instance.flip_flop_instance[22].in ),
    .RESET_B(_009_),
    .Q(\FLSR_instance.flip_flop_instance[22].out ));
 sky130_fd_sc_hd__dfrtp_1 _412_ (.CLK(net21),
    .D(\FLSR_instance.flip_flop_instance[21].in ),
    .RESET_B(_010_),
    .Q(\FLSR_instance.flip_flop_instance[21].out ));
 sky130_fd_sc_hd__dfrtp_1 _413_ (.CLK(net21),
    .D(\FLSR_instance.flip_flop_instance[20].in ),
    .RESET_B(_011_),
    .Q(\FLSR_instance.flip_flop_instance[20].out ));
 sky130_fd_sc_hd__dfrtp_1 _414_ (.CLK(net21),
    .D(\FLSR_instance.flip_flop_instance[19].in ),
    .RESET_B(_012_),
    .Q(\FLSR_instance.flip_flop_instance[19].out ));
 sky130_fd_sc_hd__dfrtp_1 _415_ (.CLK(net21),
    .D(\FLSR_instance.flip_flop_instance[18].in ),
    .RESET_B(_013_),
    .Q(\FLSR_instance.flip_flop_instance[18].out ));
 sky130_fd_sc_hd__dfrtp_1 _416_ (.CLK(net21),
    .D(\FLSR_instance.flip_flop_instance[17].in ),
    .RESET_B(_014_),
    .Q(\FLSR_instance.flip_flop_instance[17].out ));
 sky130_fd_sc_hd__dfrtp_1 _417_ (.CLK(net22),
    .D(\FLSR_instance.flip_flop_instance[16].in ),
    .RESET_B(_015_),
    .Q(\FLSR_instance.flip_flop_instance[16].out ));
 sky130_fd_sc_hd__dfrtp_1 _418_ (.CLK(net22),
    .D(\FLSR_instance.flip_flop_instance[15].in ),
    .RESET_B(_016_),
    .Q(\FLSR_instance.flip_flop_instance[15].out ));
 sky130_fd_sc_hd__dfrtp_1 _419_ (.CLK(net22),
    .D(\FLSR_instance.flip_flop_instance[14].in ),
    .RESET_B(_017_),
    .Q(\FLSR_instance.flip_flop_instance[14].out ));
 sky130_fd_sc_hd__dfrtp_1 _420_ (.CLK(net25),
    .D(\FLSR_instance.flip_flop_instance[13].in ),
    .RESET_B(_018_),
    .Q(\FLSR_instance.flip_flop_instance[13].out ));
 sky130_fd_sc_hd__dfrtp_1 _421_ (.CLK(net25),
    .D(\FLSR_instance.flip_flop_instance[12].in ),
    .RESET_B(_019_),
    .Q(\FLSR_instance.flip_flop_instance[12].out ));
 sky130_fd_sc_hd__dfrtp_1 _422_ (.CLK(net26),
    .D(\FLSR_instance.flip_flop_instance[11].in ),
    .RESET_B(_020_),
    .Q(\FLSR_instance.flip_flop_instance[11].out ));
 sky130_fd_sc_hd__dfrtp_1 _423_ (.CLK(net26),
    .D(\FLSR_instance.flip_flop_instance[10].in ),
    .RESET_B(_021_),
    .Q(\FLSR_instance.flip_flop_instance[10].out ));
 sky130_fd_sc_hd__dfrtp_1 _424_ (.CLK(net26),
    .D(\FLSR_instance.flip_flop_instance[9].in ),
    .RESET_B(_022_),
    .Q(\FLSR_instance.flip_flop_instance[9].out ));
 sky130_fd_sc_hd__dfrtp_1 _425_ (.CLK(net26),
    .D(\FLSR_instance.flip_flop_instance[8].in ),
    .RESET_B(_023_),
    .Q(\FLSR_instance.flip_flop_instance[8].out ));
 sky130_fd_sc_hd__dfrtp_1 _426_ (.CLK(net26),
    .D(\FLSR_instance.flip_flop_instance[7].in ),
    .RESET_B(_024_),
    .Q(\FLSR_instance.flip_flop_instance[7].out ));
 sky130_fd_sc_hd__dfrtp_1 _427_ (.CLK(net23),
    .D(\FLSR_instance.flip_flop_instance[6].in ),
    .RESET_B(_025_),
    .Q(\FLSR_instance.flip_flop_instance[6].out ));
 sky130_fd_sc_hd__dfrtp_1 _428_ (.CLK(net24),
    .D(\FLSR_instance.flip_flop_instance[5].in ),
    .RESET_B(_026_),
    .Q(\FLSR_instance.flip_flop_instance[5].out ));
 sky130_fd_sc_hd__dfrtp_1 _429_ (.CLK(net24),
    .D(\FLSR_instance.flip_flop_instance[4].in ),
    .RESET_B(_027_),
    .Q(\FLSR_instance.flip_flop_instance[4].out ));
 sky130_fd_sc_hd__dfrtp_1 _430_ (.CLK(net24),
    .D(\FLSR_instance.flip_flop_instance[3].in ),
    .RESET_B(_028_),
    .Q(\FLSR_instance.flip_flop_instance[3].out ));
 sky130_fd_sc_hd__dfrtp_1 _431_ (.CLK(net24),
    .D(\FLSR_instance.flip_flop_instance[2].in ),
    .RESET_B(_029_),
    .Q(\FLSR_instance.flip_flop_instance[2].out ));
 sky130_fd_sc_hd__dfrtp_1 _432_ (.CLK(net23),
    .D(\FLSR_instance.flip_flop_instance[1].in ),
    .RESET_B(_030_),
    .Q(\FLSR_instance.flip_flop_instance[1].out ));
 sky130_fd_sc_hd__dfrtp_1 _433_ (.CLK(net23),
    .D(\FLSR_instance.flip_flop_instance[0].in ),
    .RESET_B(_031_),
    .Q(\FLSR_instance.flip_flop_instance[0].out ));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net27),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 fanout20 (.A(net27),
    .X(net20));
 sky130_fd_sc_hd__buf_2 fanout21 (.A(net27),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(net27),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net27),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(net27),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(net27),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net1),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(i_clk),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(i_wb_data[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(i_wb_data[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(i_wb_data[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(i_wb_data[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(i_wb_data[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(i_wb_stb),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(i_wb_we),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(i_reset),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(i_wb_addr[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(i_wb_addr[1]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(i_wb_addr[2]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(i_wb_cyc),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(i_wb_data[0]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(i_wb_data[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(i_wb_data[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(o_wb_ack));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(o_wb_data));
 sky130_fd_sc_hd__conb_1 wb_lfsr_28 (.LO(net28));
 assign o_wb_stall = net28;
endmodule

