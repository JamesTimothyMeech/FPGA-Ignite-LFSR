magic
tech sky130A
magscale 1 2
timestamp 1692995760
<< viali >>
rect 1593 17289 1627 17323
rect 5181 17289 5215 17323
rect 5733 17289 5767 17323
rect 3433 17221 3467 17255
rect 7941 17221 7975 17255
rect 11805 17221 11839 17255
rect 15945 17221 15979 17255
rect 1501 17153 1535 17187
rect 4057 17153 4091 17187
rect 5641 17153 5675 17187
rect 9321 17153 9355 17187
rect 15577 17153 15611 17187
rect 3801 17085 3835 17119
rect 5917 17085 5951 17119
rect 9413 17085 9447 17119
rect 9505 17085 9539 17119
rect 3525 16949 3559 16983
rect 5273 16949 5307 16983
rect 8033 16949 8067 16983
rect 8953 16949 8987 16983
rect 11897 16949 11931 16983
rect 15761 16949 15795 16983
rect 16037 16949 16071 16983
rect 3893 16745 3927 16779
rect 6929 16745 6963 16779
rect 8769 16745 8803 16779
rect 1685 16609 1719 16643
rect 4813 16609 4847 16643
rect 5181 16609 5215 16643
rect 5457 16609 5491 16643
rect 7021 16609 7055 16643
rect 9045 16609 9079 16643
rect 1409 16541 1443 16575
rect 4077 16541 4111 16575
rect 4629 16541 4663 16575
rect 1952 16473 1986 16507
rect 7297 16473 7331 16507
rect 9312 16473 9346 16507
rect 1593 16405 1627 16439
rect 3065 16405 3099 16439
rect 4261 16405 4295 16439
rect 4721 16405 4755 16439
rect 10425 16405 10459 16439
rect 2145 16201 2179 16235
rect 2605 16201 2639 16235
rect 6469 16201 6503 16235
rect 7021 16201 7055 16235
rect 7481 16201 7515 16235
rect 8401 16201 8435 16235
rect 9321 16201 9355 16235
rect 9781 16201 9815 16235
rect 11161 16201 11195 16235
rect 13277 16201 13311 16235
rect 13737 16201 13771 16235
rect 3065 16133 3099 16167
rect 3801 16133 3835 16167
rect 11805 16133 11839 16167
rect 2329 16065 2363 16099
rect 2973 16065 3007 16099
rect 3617 16065 3651 16099
rect 4445 16065 4479 16099
rect 6653 16065 6687 16099
rect 6929 16065 6963 16099
rect 7665 16065 7699 16099
rect 8309 16065 8343 16099
rect 9965 16065 9999 16099
rect 11345 16065 11379 16099
rect 3249 15997 3283 16031
rect 3433 15997 3467 16031
rect 4721 15997 4755 16031
rect 9413 15997 9447 16031
rect 9597 15997 9631 16031
rect 11529 15997 11563 16031
rect 13829 15997 13863 16031
rect 13921 15997 13955 16031
rect 8953 15929 8987 15963
rect 6193 15861 6227 15895
rect 13369 15861 13403 15895
rect 5273 15657 5307 15691
rect 6285 15657 6319 15691
rect 9413 15657 9447 15691
rect 12265 15657 12299 15691
rect 5181 15589 5215 15623
rect 9045 15521 9079 15555
rect 4905 15453 4939 15487
rect 4997 15453 5031 15487
rect 5457 15453 5491 15487
rect 6193 15453 6227 15487
rect 9229 15453 9263 15487
rect 12173 15453 12207 15487
rect 13001 15453 13035 15487
rect 14105 15453 14139 15487
rect 9781 15317 9815 15351
rect 12817 15317 12851 15351
rect 14197 15317 14231 15351
rect 2789 15113 2823 15147
rect 7389 15113 7423 15147
rect 11345 15113 11379 15147
rect 11897 15113 11931 15147
rect 13185 15045 13219 15079
rect 1676 14977 1710 15011
rect 7757 14977 7791 15011
rect 8309 14977 8343 15011
rect 9597 14977 9631 15011
rect 12909 14977 12943 15011
rect 1409 14909 1443 14943
rect 7849 14909 7883 14943
rect 8033 14909 8067 14943
rect 9873 14909 9907 14943
rect 11989 14909 12023 14943
rect 12081 14909 12115 14943
rect 11529 14841 11563 14875
rect 8401 14773 8435 14807
rect 14657 14773 14691 14807
rect 1685 14569 1719 14603
rect 7389 14569 7423 14603
rect 9781 14569 9815 14603
rect 10701 14569 10735 14603
rect 13185 14569 13219 14603
rect 5181 14501 5215 14535
rect 5273 14501 5307 14535
rect 8953 14501 8987 14535
rect 2605 14433 2639 14467
rect 3801 14433 3835 14467
rect 5917 14433 5951 14467
rect 9597 14433 9631 14467
rect 11805 14433 11839 14467
rect 14657 14433 14691 14467
rect 1869 14365 1903 14399
rect 2329 14365 2363 14399
rect 3157 14365 3191 14399
rect 3341 14365 3375 14399
rect 3433 14365 3467 14399
rect 5457 14365 5491 14399
rect 5641 14365 5675 14399
rect 7481 14365 7515 14399
rect 8033 14365 8067 14399
rect 9413 14365 9447 14399
rect 9965 14365 9999 14399
rect 10609 14365 10643 14399
rect 14473 14365 14507 14399
rect 4046 14297 4080 14331
rect 7573 14297 7607 14331
rect 9321 14297 9355 14331
rect 12072 14297 12106 14331
rect 1961 14229 1995 14263
rect 2421 14229 2455 14263
rect 2973 14229 3007 14263
rect 3617 14229 3651 14263
rect 7849 14229 7883 14263
rect 14105 14229 14139 14263
rect 14565 14229 14599 14263
rect 1869 14025 1903 14059
rect 2237 14025 2271 14059
rect 2697 14025 2731 14059
rect 3433 14025 3467 14059
rect 3893 14025 3927 14059
rect 4353 14025 4387 14059
rect 4813 14025 4847 14059
rect 5733 14025 5767 14059
rect 8861 14025 8895 14059
rect 9321 14025 9355 14059
rect 9965 14025 9999 14059
rect 12357 14025 12391 14059
rect 16221 14025 16255 14059
rect 3801 13957 3835 13991
rect 7748 13957 7782 13991
rect 12081 13957 12115 13991
rect 14473 13957 14507 13991
rect 2053 13889 2087 13923
rect 2605 13889 2639 13923
rect 4721 13889 4755 13923
rect 5365 13889 5399 13923
rect 7481 13889 7515 13923
rect 9045 13889 9079 13923
rect 9137 13889 9171 13923
rect 10333 13889 10367 13923
rect 10425 13889 10459 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 12173 13889 12207 13923
rect 13165 13889 13199 13923
rect 14381 13889 14415 13923
rect 14841 13889 14875 13923
rect 16037 13889 16071 13923
rect 2881 13821 2915 13855
rect 4077 13821 4111 13855
rect 4997 13821 5031 13855
rect 5273 13821 5307 13855
rect 10517 13821 10551 13855
rect 12909 13821 12943 13855
rect 14657 13753 14691 13787
rect 14289 13685 14323 13719
rect 5089 13481 5123 13515
rect 10701 13481 10735 13515
rect 12173 13481 12207 13515
rect 12909 13481 12943 13515
rect 3341 13345 3375 13379
rect 4721 13345 4755 13379
rect 8953 13345 8987 13379
rect 14105 13345 14139 13379
rect 14381 13345 14415 13379
rect 4813 13277 4847 13311
rect 8125 13277 8159 13311
rect 10793 13277 10827 13311
rect 12357 13277 12391 13311
rect 12725 13277 12759 13311
rect 9229 13209 9263 13243
rect 11060 13209 11094 13243
rect 12541 13209 12575 13243
rect 12633 13209 12667 13243
rect 2697 13141 2731 13175
rect 3065 13141 3099 13175
rect 3157 13141 3191 13175
rect 7941 13141 7975 13175
rect 15853 13141 15887 13175
rect 2605 12937 2639 12971
rect 4629 12937 4663 12971
rect 5825 12937 5859 12971
rect 8769 12937 8803 12971
rect 9045 12937 9079 12971
rect 9505 12937 9539 12971
rect 11345 12937 11379 12971
rect 13277 12937 13311 12971
rect 3157 12869 3191 12903
rect 8585 12869 8619 12903
rect 10517 12869 10551 12903
rect 10977 12869 11011 12903
rect 11069 12869 11103 12903
rect 12173 12869 12207 12903
rect 12265 12869 12299 12903
rect 13369 12869 13403 12903
rect 1501 12801 1535 12835
rect 2329 12801 2363 12835
rect 2789 12801 2823 12835
rect 2881 12801 2915 12835
rect 8953 12801 8987 12835
rect 9413 12801 9447 12835
rect 10241 12801 10275 12835
rect 10793 12801 10827 12835
rect 11161 12801 11195 12835
rect 11989 12801 12023 12835
rect 12357 12801 12391 12835
rect 14013 12801 14047 12835
rect 5917 12733 5951 12767
rect 6101 12733 6135 12767
rect 6377 12733 6411 12767
rect 6653 12733 6687 12767
rect 13553 12733 13587 12767
rect 13737 12733 13771 12767
rect 2421 12665 2455 12699
rect 8217 12665 8251 12699
rect 1593 12597 1627 12631
rect 5457 12597 5491 12631
rect 8125 12597 8159 12631
rect 8585 12597 8619 12631
rect 12541 12597 12575 12631
rect 12909 12597 12943 12631
rect 3157 12393 3191 12427
rect 3985 12393 4019 12427
rect 5181 12393 5215 12427
rect 5733 12393 5767 12427
rect 6929 12393 6963 12427
rect 7297 12393 7331 12427
rect 12173 12393 12207 12427
rect 13645 12393 13679 12427
rect 1409 12257 1443 12291
rect 1685 12257 1719 12291
rect 4905 12257 4939 12291
rect 7941 12257 7975 12291
rect 9229 12257 9263 12291
rect 3893 12189 3927 12223
rect 4813 12189 4847 12223
rect 5917 12189 5951 12223
rect 6837 12189 6871 12223
rect 10793 12189 10827 12223
rect 12265 12189 12299 12223
rect 12532 12189 12566 12223
rect 14289 12189 14323 12223
rect 9474 12121 9508 12155
rect 11060 12121 11094 12155
rect 7665 12053 7699 12087
rect 7757 12053 7791 12087
rect 10609 12053 10643 12087
rect 14105 12053 14139 12087
rect 9229 11849 9263 11883
rect 12081 11849 12115 11883
rect 11713 11781 11747 11815
rect 11805 11781 11839 11815
rect 14013 11781 14047 11815
rect 2605 11713 2639 11747
rect 6561 11713 6595 11747
rect 6817 11713 6851 11747
rect 9413 11713 9447 11747
rect 11529 11713 11563 11747
rect 11897 11713 11931 11747
rect 13737 11713 13771 11747
rect 2421 11509 2455 11543
rect 7941 11509 7975 11543
rect 15485 11509 15519 11543
rect 3341 11305 3375 11339
rect 6009 11305 6043 11339
rect 8585 11305 8619 11339
rect 9137 11305 9171 11339
rect 15853 11305 15887 11339
rect 6101 11237 6135 11271
rect 8769 11237 8803 11271
rect 12173 11237 12207 11271
rect 13645 11237 13679 11271
rect 14381 11237 14415 11271
rect 15761 11237 15795 11271
rect 3801 11169 3835 11203
rect 6745 11169 6779 11203
rect 7665 11169 7699 11203
rect 9689 11169 9723 11203
rect 10977 11169 11011 11203
rect 14841 11169 14875 11203
rect 14933 11169 14967 11203
rect 1869 11101 1903 11135
rect 1961 11101 1995 11135
rect 2228 11101 2262 11135
rect 3985 11101 4019 11135
rect 4629 11101 4663 11135
rect 6469 11101 6503 11135
rect 7389 11101 7423 11135
rect 9505 11101 9539 11135
rect 10701 11101 10735 11135
rect 11621 11101 11655 11135
rect 11805 11101 11839 11135
rect 11989 11101 12023 11135
rect 12265 11101 12299 11135
rect 12521 11101 12555 11135
rect 14749 11101 14783 11135
rect 4874 11033 4908 11067
rect 6561 11033 6595 11067
rect 8401 11033 8435 11067
rect 9597 11033 9631 11067
rect 11897 11033 11931 11067
rect 15393 11033 15427 11067
rect 1685 10965 1719 10999
rect 4169 10965 4203 10999
rect 7021 10965 7055 10999
rect 7481 10965 7515 10999
rect 8601 10965 8635 10999
rect 2881 10761 2915 10795
rect 3249 10761 3283 10795
rect 4997 10761 5031 10795
rect 5825 10761 5859 10795
rect 6837 10761 6871 10795
rect 7481 10761 7515 10795
rect 8953 10761 8987 10795
rect 9597 10761 9631 10795
rect 10977 10761 11011 10795
rect 11713 10761 11747 10795
rect 14933 10761 14967 10795
rect 1676 10693 1710 10727
rect 10517 10693 10551 10727
rect 1409 10625 1443 10659
rect 3341 10625 3375 10659
rect 4077 10625 4111 10659
rect 5181 10625 5215 10659
rect 5641 10625 5675 10659
rect 7021 10625 7055 10659
rect 7297 10625 7331 10659
rect 8217 10625 8251 10659
rect 8769 10625 8803 10659
rect 8861 10625 8895 10659
rect 9413 10625 9447 10659
rect 9597 10625 9631 10659
rect 11069 10625 11103 10659
rect 11253 10625 11287 10659
rect 11529 10625 11563 10659
rect 14473 10625 14507 10659
rect 14841 10625 14875 10659
rect 15301 10625 15335 10659
rect 3525 10557 3559 10591
rect 4353 10557 4387 10591
rect 5457 10557 5491 10591
rect 7113 10557 7147 10591
rect 8033 10557 8067 10591
rect 8401 10557 8435 10591
rect 9229 10557 9263 10591
rect 9781 10557 9815 10591
rect 10517 10489 10551 10523
rect 2789 10421 2823 10455
rect 8493 10421 8527 10455
rect 9137 10421 9171 10455
rect 14657 10421 14691 10455
rect 15117 10421 15151 10455
rect 5549 10217 5583 10251
rect 9689 10217 9723 10251
rect 9965 10217 9999 10251
rect 11437 10217 11471 10251
rect 13921 10217 13955 10251
rect 3801 10081 3835 10115
rect 6377 10081 6411 10115
rect 9689 10081 9723 10115
rect 12541 10081 12575 10115
rect 14749 10081 14783 10115
rect 3617 10013 3651 10047
rect 5733 10013 5767 10047
rect 9597 10013 9631 10047
rect 11253 10013 11287 10047
rect 11897 10013 11931 10047
rect 12081 10013 12115 10047
rect 12173 10013 12207 10047
rect 12265 10013 12299 10047
rect 14473 10013 14507 10047
rect 4077 9945 4111 9979
rect 6644 9945 6678 9979
rect 9137 9945 9171 9979
rect 12786 9945 12820 9979
rect 3433 9877 3467 9911
rect 6009 9877 6043 9911
rect 7757 9877 7791 9911
rect 9413 9877 9447 9911
rect 12449 9877 12483 9911
rect 16221 9877 16255 9911
rect 3525 9673 3559 9707
rect 4537 9673 4571 9707
rect 6653 9673 6687 9707
rect 6929 9673 6963 9707
rect 14565 9673 14599 9707
rect 15393 9673 15427 9707
rect 7849 9605 7883 9639
rect 7941 9605 7975 9639
rect 8401 9605 8435 9639
rect 10977 9605 11011 9639
rect 14657 9605 14691 9639
rect 1409 9537 1443 9571
rect 1676 9537 1710 9571
rect 3893 9537 3927 9571
rect 4445 9537 4479 9571
rect 6469 9537 6503 9571
rect 7113 9537 7147 9571
rect 8309 9537 8343 9571
rect 8493 9537 8527 9571
rect 8953 9537 8987 9571
rect 10149 9537 10183 9571
rect 10793 9537 10827 9571
rect 11069 9537 11103 9571
rect 11161 9537 11195 9571
rect 11785 9537 11819 9571
rect 15209 9537 15243 9571
rect 15301 9537 15335 9571
rect 16313 9537 16347 9571
rect 3985 9469 4019 9503
rect 4077 9469 4111 9503
rect 8125 9469 8159 9503
rect 9229 9469 9263 9503
rect 11529 9469 11563 9503
rect 14841 9469 14875 9503
rect 2789 9401 2823 9435
rect 7481 9401 7515 9435
rect 11345 9401 11379 9435
rect 12909 9401 12943 9435
rect 14197 9401 14231 9435
rect 9321 9333 9355 9367
rect 9505 9333 9539 9367
rect 10241 9333 10275 9367
rect 15025 9333 15059 9367
rect 1593 9129 1627 9163
rect 7941 9129 7975 9163
rect 8769 9129 8803 9163
rect 10241 9129 10275 9163
rect 11161 9129 11195 9163
rect 11437 9129 11471 9163
rect 11713 9129 11747 9163
rect 10701 9061 10735 9095
rect 10885 9061 10919 9095
rect 2513 8993 2547 9027
rect 5457 8993 5491 9027
rect 8953 8993 8987 9027
rect 10425 8993 10459 9027
rect 13093 8993 13127 9027
rect 13277 8993 13311 9027
rect 14381 8993 14415 9027
rect 1777 8925 1811 8959
rect 2237 8925 2271 8959
rect 3893 8925 3927 8959
rect 5365 8925 5399 8959
rect 5641 8925 5675 8959
rect 7849 8925 7883 8959
rect 8217 8925 8251 8959
rect 8585 8925 8619 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 9781 8925 9815 8959
rect 9873 8925 9907 8959
rect 10977 8925 11011 8959
rect 14105 8925 14139 8959
rect 15945 8925 15979 8959
rect 11529 8857 11563 8891
rect 11729 8857 11763 8891
rect 13001 8857 13035 8891
rect 16037 8857 16071 8891
rect 1869 8789 1903 8823
rect 2329 8789 2363 8823
rect 3985 8789 4019 8823
rect 5181 8789 5215 8823
rect 5825 8789 5859 8823
rect 8401 8789 8435 8823
rect 11897 8789 11931 8823
rect 12633 8789 12667 8823
rect 15853 8789 15887 8823
rect 2421 8585 2455 8619
rect 4353 8585 4387 8619
rect 2881 8517 2915 8551
rect 5080 8517 5114 8551
rect 1409 8449 1443 8483
rect 2237 8449 2271 8483
rect 2605 8449 2639 8483
rect 7021 8449 7055 8483
rect 8493 8449 8527 8483
rect 8677 8449 8711 8483
rect 8861 8449 8895 8483
rect 9321 8449 9355 8483
rect 9413 8449 9447 8483
rect 10149 8449 10183 8483
rect 10701 8449 10735 8483
rect 11069 8449 11103 8483
rect 12909 8449 12943 8483
rect 2053 8381 2087 8415
rect 4813 8381 4847 8415
rect 1593 8313 1627 8347
rect 11069 8313 11103 8347
rect 6193 8245 6227 8279
rect 6837 8245 6871 8279
rect 9781 8245 9815 8279
rect 12725 8245 12759 8279
rect 2973 8041 3007 8075
rect 5365 8041 5399 8075
rect 9321 8041 9355 8075
rect 4445 7905 4479 7939
rect 5825 7905 5859 7939
rect 6009 7905 6043 7939
rect 7941 7905 7975 7939
rect 12449 7905 12483 7939
rect 14749 7905 14783 7939
rect 3157 7837 3191 7871
rect 5733 7837 5767 7871
rect 6469 7837 6503 7871
rect 6725 7837 6759 7871
rect 8125 7837 8159 7871
rect 8953 7837 8987 7871
rect 9597 7837 9631 7871
rect 9689 7837 9723 7871
rect 10057 7837 10091 7871
rect 10885 7837 10919 7871
rect 11529 7837 11563 7871
rect 11897 7837 11931 7871
rect 12173 7837 12207 7871
rect 14565 7837 14599 7871
rect 4261 7769 4295 7803
rect 9330 7769 9364 7803
rect 9873 7769 9907 7803
rect 9965 7769 9999 7803
rect 11713 7769 11747 7803
rect 11805 7769 11839 7803
rect 14473 7769 14507 7803
rect 3801 7701 3835 7735
rect 4169 7701 4203 7735
rect 7849 7701 7883 7735
rect 8309 7701 8343 7735
rect 10241 7701 10275 7735
rect 11069 7701 11103 7735
rect 12081 7701 12115 7735
rect 13921 7701 13955 7735
rect 14105 7701 14139 7735
rect 2789 7497 2823 7531
rect 4905 7497 4939 7531
rect 5733 7497 5767 7531
rect 7021 7497 7055 7531
rect 7389 7497 7423 7531
rect 7481 7497 7515 7531
rect 13369 7497 13403 7531
rect 13737 7497 13771 7531
rect 5089 7429 5123 7463
rect 8760 7429 8794 7463
rect 12234 7429 12268 7463
rect 1409 7361 1443 7395
rect 1676 7361 1710 7395
rect 4997 7361 5031 7395
rect 5641 7361 5675 7395
rect 8493 7361 8527 7395
rect 9965 7361 9999 7395
rect 10232 7361 10266 7395
rect 11989 7361 12023 7395
rect 13645 7361 13679 7395
rect 14197 7361 14231 7395
rect 15025 7361 15059 7395
rect 3157 7293 3191 7327
rect 3433 7293 3467 7327
rect 5917 7293 5951 7327
rect 7665 7293 7699 7327
rect 5273 7157 5307 7191
rect 9873 7157 9907 7191
rect 11345 7157 11379 7191
rect 14013 7157 14047 7191
rect 15117 7157 15151 7191
rect 1685 6953 1719 6987
rect 3893 6953 3927 6987
rect 11069 6953 11103 6987
rect 14362 6953 14396 6987
rect 2513 6817 2547 6851
rect 7389 6817 7423 6851
rect 7481 6817 7515 6851
rect 9505 6817 9539 6851
rect 13921 6817 13955 6851
rect 14105 6817 14139 6851
rect 1869 6749 1903 6783
rect 2329 6749 2363 6783
rect 2789 6749 2823 6783
rect 2973 6749 3007 6783
rect 4077 6749 4111 6783
rect 9413 6749 9447 6783
rect 10517 6749 10551 6783
rect 10885 6749 10919 6783
rect 5917 6681 5951 6715
rect 10701 6681 10735 6715
rect 10793 6681 10827 6715
rect 13737 6681 13771 6715
rect 1961 6613 1995 6647
rect 2421 6613 2455 6647
rect 3157 6613 3191 6647
rect 6009 6613 6043 6647
rect 6929 6613 6963 6647
rect 7297 6613 7331 6647
rect 8953 6613 8987 6647
rect 9321 6613 9355 6647
rect 15853 6613 15887 6647
rect 8125 6409 8159 6443
rect 12265 6409 12299 6443
rect 14657 6409 14691 6443
rect 12602 6341 12636 6375
rect 3433 6273 3467 6307
rect 4261 6273 4295 6307
rect 6377 6273 6411 6307
rect 8861 6273 8895 6307
rect 11713 6273 11747 6307
rect 11897 6273 11931 6307
rect 11989 6273 12023 6307
rect 12081 6273 12115 6307
rect 4537 6205 4571 6239
rect 6653 6205 6687 6239
rect 12357 6205 12391 6239
rect 14749 6205 14783 6239
rect 14933 6205 14967 6239
rect 6009 6137 6043 6171
rect 13737 6137 13771 6171
rect 3249 6069 3283 6103
rect 8677 6069 8711 6103
rect 14289 6069 14323 6103
rect 4813 5865 4847 5899
rect 5365 5865 5399 5899
rect 6193 5865 6227 5899
rect 6837 5865 6871 5899
rect 9137 5865 9171 5899
rect 16129 5865 16163 5899
rect 8769 5797 8803 5831
rect 2697 5729 2731 5763
rect 7021 5729 7055 5763
rect 7297 5729 7331 5763
rect 9689 5729 9723 5763
rect 10149 5729 10183 5763
rect 12449 5729 12483 5763
rect 12541 5729 12575 5763
rect 2881 5661 2915 5695
rect 3893 5661 3927 5695
rect 4997 5661 5031 5695
rect 5273 5661 5307 5695
rect 6377 5661 6411 5695
rect 6745 5661 6779 5695
rect 12817 5661 12851 5695
rect 14565 5661 14599 5695
rect 16313 5661 16347 5695
rect 9505 5593 9539 5627
rect 10425 5593 10459 5627
rect 12909 5593 12943 5627
rect 3065 5525 3099 5559
rect 3985 5525 4019 5559
rect 9597 5525 9631 5559
rect 11897 5525 11931 5559
rect 11989 5525 12023 5559
rect 12357 5525 12391 5559
rect 14381 5525 14415 5559
rect 1869 5321 1903 5355
rect 2329 5321 2363 5355
rect 7941 5321 7975 5355
rect 10057 5321 10091 5355
rect 10517 5321 10551 5355
rect 12173 5321 12207 5355
rect 2237 5253 2271 5287
rect 2973 5253 3007 5287
rect 12510 5253 12544 5287
rect 14473 5253 14507 5287
rect 16129 5253 16163 5287
rect 1777 5185 1811 5219
rect 2697 5185 2731 5219
rect 5457 5185 5491 5219
rect 7849 5185 7883 5219
rect 8677 5185 8711 5219
rect 8944 5185 8978 5219
rect 10701 5185 10735 5219
rect 11621 5185 11655 5219
rect 11805 5185 11839 5219
rect 11897 5185 11931 5219
rect 11989 5185 12023 5219
rect 12265 5185 12299 5219
rect 14197 5185 14231 5219
rect 16037 5185 16071 5219
rect 2513 5117 2547 5151
rect 1593 4981 1627 5015
rect 4445 4981 4479 5015
rect 5273 4981 5307 5015
rect 13645 4981 13679 5015
rect 15945 4981 15979 5015
rect 4721 4777 4755 4811
rect 9781 4777 9815 4811
rect 2789 4709 2823 4743
rect 5365 4641 5399 4675
rect 5825 4641 5859 4675
rect 14565 4641 14599 4675
rect 14749 4641 14783 4675
rect 1409 4573 1443 4607
rect 1676 4573 1710 4607
rect 3985 4573 4019 4607
rect 4353 4573 4387 4607
rect 5089 4573 5123 4607
rect 5549 4573 5583 4607
rect 7389 4573 7423 4607
rect 7665 4573 7699 4607
rect 9229 4573 9263 4607
rect 9413 4573 9447 4607
rect 9597 4573 9631 4607
rect 10333 4573 10367 4607
rect 13921 4573 13955 4607
rect 14473 4573 14507 4607
rect 7481 4505 7515 4539
rect 9505 4505 9539 4539
rect 3801 4437 3835 4471
rect 4445 4437 4479 4471
rect 5181 4437 5215 4471
rect 7297 4437 7331 4471
rect 7757 4437 7791 4471
rect 10149 4437 10183 4471
rect 13737 4437 13771 4471
rect 14105 4437 14139 4471
rect 5181 4233 5215 4267
rect 5641 4233 5675 4267
rect 8493 4233 8527 4267
rect 13093 4233 13127 4267
rect 15485 4233 15519 4267
rect 1501 4165 1535 4199
rect 3709 4165 3743 4199
rect 9873 4165 9907 4199
rect 1685 4097 1719 4131
rect 6653 4097 6687 4131
rect 11529 4097 11563 4131
rect 11621 4097 11655 4131
rect 12541 4097 12575 4131
rect 13737 4097 13771 4131
rect 15577 4097 15611 4131
rect 15669 4097 15703 4131
rect 3433 4029 3467 4063
rect 5733 4029 5767 4063
rect 5825 4029 5859 4063
rect 6745 4029 6779 4063
rect 7021 4029 7055 4063
rect 9597 4029 9631 4063
rect 11345 4029 11379 4063
rect 13185 4029 13219 4063
rect 13369 4029 13403 4063
rect 14013 4029 14047 4063
rect 6469 3961 6503 3995
rect 12725 3961 12759 3995
rect 5273 3893 5307 3927
rect 12357 3893 12391 3927
rect 3801 3689 3835 3723
rect 7021 3689 7055 3723
rect 10333 3689 10367 3723
rect 14657 3689 14691 3723
rect 14289 3621 14323 3655
rect 4445 3553 4479 3587
rect 7573 3553 7607 3587
rect 10977 3553 11011 3587
rect 11897 3553 11931 3587
rect 12173 3553 12207 3587
rect 2973 3485 3007 3519
rect 4169 3485 4203 3519
rect 4905 3485 4939 3519
rect 5181 3485 5215 3519
rect 5273 3485 5307 3519
rect 7389 3485 7423 3519
rect 13737 3485 13771 3519
rect 14105 3485 14139 3519
rect 14473 3485 14507 3519
rect 13829 3417 13863 3451
rect 2789 3349 2823 3383
rect 4261 3349 4295 3383
rect 4721 3349 4755 3383
rect 5457 3349 5491 3383
rect 7481 3349 7515 3383
rect 10701 3349 10735 3383
rect 10793 3349 10827 3383
rect 13645 3349 13679 3383
rect 3801 3145 3835 3179
rect 5825 3145 5859 3179
rect 7849 3145 7883 3179
rect 8309 3145 8343 3179
rect 13369 3145 13403 3179
rect 2688 3077 2722 3111
rect 4701 3077 4735 3111
rect 8401 3077 8435 3111
rect 9137 3077 9171 3111
rect 2421 3009 2455 3043
rect 3893 3009 3927 3043
rect 4077 3009 4111 3043
rect 4445 3009 4479 3043
rect 6469 3009 6503 3043
rect 6736 3009 6770 3043
rect 8953 3009 8987 3043
rect 9781 3009 9815 3043
rect 10048 3009 10082 3043
rect 11989 3009 12023 3043
rect 12256 3009 12290 3043
rect 8493 2941 8527 2975
rect 8769 2941 8803 2975
rect 4261 2805 4295 2839
rect 7941 2805 7975 2839
rect 11161 2805 11195 2839
rect 2881 2601 2915 2635
rect 4905 2601 4939 2635
rect 6745 2601 6779 2635
rect 7021 2601 7055 2635
rect 8033 2601 8067 2635
rect 10517 2601 10551 2635
rect 12357 2601 12391 2635
rect 12633 2601 12667 2635
rect 16129 2601 16163 2635
rect 1593 2533 1627 2567
rect 15853 2533 15887 2567
rect 3525 2465 3559 2499
rect 5457 2465 5491 2499
rect 1409 2397 1443 2431
rect 3341 2397 3375 2431
rect 5365 2397 5399 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 7849 2397 7883 2431
rect 9965 2397 9999 2431
rect 10333 2397 10367 2431
rect 11805 2397 11839 2431
rect 12173 2397 12207 2431
rect 12449 2397 12483 2431
rect 16313 2397 16347 2431
rect 3249 2329 3283 2363
rect 4077 2329 4111 2363
rect 5273 2329 5307 2363
rect 10149 2329 10183 2363
rect 10241 2329 10275 2363
rect 11989 2329 12023 2363
rect 12081 2329 12115 2363
rect 15669 2329 15703 2363
rect 4169 2261 4203 2295
<< metal1 >>
rect 1104 17434 16811 17456
rect 1104 17382 4836 17434
rect 4888 17382 4900 17434
rect 4952 17382 4964 17434
rect 5016 17382 5028 17434
rect 5080 17382 5092 17434
rect 5144 17382 8723 17434
rect 8775 17382 8787 17434
rect 8839 17382 8851 17434
rect 8903 17382 8915 17434
rect 8967 17382 8979 17434
rect 9031 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 16497 17434
rect 16549 17382 16561 17434
rect 16613 17382 16625 17434
rect 16677 17382 16689 17434
rect 16741 17382 16753 17434
rect 16805 17382 16811 17434
rect 1104 17360 16811 17382
rect 14 17280 20 17332
rect 72 17320 78 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 72 17292 1593 17320
rect 72 17280 78 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 1581 17283 1639 17289
rect 4614 17280 4620 17332
rect 4672 17320 4678 17332
rect 5169 17323 5227 17329
rect 5169 17320 5181 17323
rect 4672 17292 5181 17320
rect 4672 17280 4678 17292
rect 5169 17289 5181 17292
rect 5215 17320 5227 17323
rect 5721 17323 5779 17329
rect 5721 17320 5733 17323
rect 5215 17292 5733 17320
rect 5215 17289 5227 17292
rect 5169 17283 5227 17289
rect 5721 17289 5733 17292
rect 5767 17289 5779 17323
rect 5721 17283 5779 17289
rect 15470 17280 15476 17332
rect 15528 17280 15534 17332
rect 3421 17255 3479 17261
rect 3421 17221 3433 17255
rect 3467 17252 3479 17255
rect 3602 17252 3608 17264
rect 3467 17224 3608 17252
rect 3467 17221 3479 17224
rect 3421 17215 3479 17221
rect 3602 17212 3608 17224
rect 3660 17212 3666 17264
rect 7742 17212 7748 17264
rect 7800 17252 7806 17264
rect 7929 17255 7987 17261
rect 7929 17252 7941 17255
rect 7800 17224 7941 17252
rect 7800 17212 7806 17224
rect 7929 17221 7941 17224
rect 7975 17221 7987 17255
rect 7929 17215 7987 17221
rect 11606 17212 11612 17264
rect 11664 17252 11670 17264
rect 11793 17255 11851 17261
rect 11793 17252 11805 17255
rect 11664 17224 11805 17252
rect 11664 17212 11670 17224
rect 11793 17221 11805 17224
rect 11839 17221 11851 17255
rect 11793 17215 11851 17221
rect 1486 17144 1492 17196
rect 1544 17144 1550 17196
rect 3878 17144 3884 17196
rect 3936 17184 3942 17196
rect 4045 17187 4103 17193
rect 4045 17184 4057 17187
rect 3936 17156 4057 17184
rect 3936 17144 3942 17156
rect 4045 17153 4057 17156
rect 4091 17153 4103 17187
rect 4045 17147 4103 17153
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 7098 17184 7104 17196
rect 5675 17156 7104 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 9306 17144 9312 17196
rect 9364 17144 9370 17196
rect 15488 17184 15516 17280
rect 15930 17212 15936 17264
rect 15988 17212 15994 17264
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 15488 17156 15577 17184
rect 15565 17153 15577 17156
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 3786 17076 3792 17128
rect 3844 17076 3850 17128
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17085 5963 17119
rect 5905 17079 5963 17085
rect 5920 17048 5948 17079
rect 9398 17076 9404 17128
rect 9456 17076 9462 17128
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 8294 17048 8300 17060
rect 5920 17020 8300 17048
rect 8294 17008 8300 17020
rect 8352 17048 8358 17060
rect 9508 17048 9536 17079
rect 8352 17020 9536 17048
rect 8352 17008 8358 17020
rect 10134 17008 10140 17060
rect 10192 17048 10198 17060
rect 10192 17020 16068 17048
rect 10192 17008 10198 17020
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 3513 16983 3571 16989
rect 3513 16980 3525 16983
rect 3384 16952 3525 16980
rect 3384 16940 3390 16952
rect 3513 16949 3525 16952
rect 3559 16949 3571 16983
rect 3513 16943 3571 16949
rect 5258 16940 5264 16992
rect 5316 16940 5322 16992
rect 8018 16940 8024 16992
rect 8076 16940 8082 16992
rect 8110 16940 8116 16992
rect 8168 16980 8174 16992
rect 8941 16983 8999 16989
rect 8941 16980 8953 16983
rect 8168 16952 8953 16980
rect 8168 16940 8174 16952
rect 8941 16949 8953 16952
rect 8987 16949 8999 16983
rect 8941 16943 8999 16949
rect 11882 16940 11888 16992
rect 11940 16940 11946 16992
rect 15746 16940 15752 16992
rect 15804 16940 15810 16992
rect 16040 16989 16068 17020
rect 16025 16983 16083 16989
rect 16025 16949 16037 16983
rect 16071 16949 16083 16983
rect 16025 16943 16083 16949
rect 1104 16890 16652 16912
rect 1104 16838 2893 16890
rect 2945 16838 2957 16890
rect 3009 16838 3021 16890
rect 3073 16838 3085 16890
rect 3137 16838 3149 16890
rect 3201 16838 6780 16890
rect 6832 16838 6844 16890
rect 6896 16838 6908 16890
rect 6960 16838 6972 16890
rect 7024 16838 7036 16890
rect 7088 16838 10667 16890
rect 10719 16838 10731 16890
rect 10783 16838 10795 16890
rect 10847 16838 10859 16890
rect 10911 16838 10923 16890
rect 10975 16838 14554 16890
rect 14606 16838 14618 16890
rect 14670 16838 14682 16890
rect 14734 16838 14746 16890
rect 14798 16838 14810 16890
rect 14862 16838 16652 16890
rect 1104 16816 16652 16838
rect 3234 16776 3240 16788
rect 1688 16748 3240 16776
rect 1688 16649 1716 16748
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 3878 16736 3884 16788
rect 3936 16736 3942 16788
rect 6917 16779 6975 16785
rect 5184 16748 6592 16776
rect 3786 16668 3792 16720
rect 3844 16708 3850 16720
rect 5184 16708 5212 16748
rect 3844 16680 5212 16708
rect 3844 16668 3850 16680
rect 1673 16643 1731 16649
rect 1673 16609 1685 16643
rect 1719 16609 1731 16643
rect 1673 16603 1731 16609
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 5184 16649 5212 16680
rect 4801 16643 4859 16649
rect 4801 16640 4813 16643
rect 4212 16612 4813 16640
rect 4212 16600 4218 16612
rect 4801 16609 4813 16612
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 5169 16643 5227 16649
rect 5169 16609 5181 16643
rect 5215 16609 5227 16643
rect 5169 16603 5227 16609
rect 5445 16643 5503 16649
rect 5445 16609 5457 16643
rect 5491 16640 5503 16643
rect 6454 16640 6460 16652
rect 5491 16612 6460 16640
rect 5491 16609 5503 16612
rect 5445 16603 5503 16609
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 6564 16640 6592 16748
rect 6917 16745 6929 16779
rect 6963 16776 6975 16779
rect 7098 16776 7104 16788
rect 6963 16748 7104 16776
rect 6963 16745 6975 16748
rect 6917 16739 6975 16745
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 9306 16776 9312 16788
rect 8803 16748 9312 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 7009 16643 7067 16649
rect 7009 16640 7021 16643
rect 6564 16612 7021 16640
rect 7009 16609 7021 16612
rect 7055 16609 7067 16643
rect 7009 16603 7067 16609
rect 9033 16643 9091 16649
rect 9033 16609 9045 16643
rect 9079 16640 9091 16643
rect 11054 16640 11060 16652
rect 9079 16612 9168 16640
rect 9079 16609 9091 16612
rect 9033 16603 9091 16609
rect 934 16532 940 16584
rect 992 16572 998 16584
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 992 16544 1409 16572
rect 992 16532 998 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 4111 16544 4292 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 1940 16507 1998 16513
rect 1940 16473 1952 16507
rect 1986 16504 1998 16507
rect 2130 16504 2136 16516
rect 1986 16476 2136 16504
rect 1986 16473 1998 16476
rect 1940 16467 1998 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16436 1639 16439
rect 2682 16436 2688 16448
rect 1627 16408 2688 16436
rect 1627 16405 1639 16408
rect 1581 16399 1639 16405
rect 2682 16396 2688 16408
rect 2740 16396 2746 16448
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 4264 16445 4292 16544
rect 4614 16532 4620 16584
rect 4672 16532 4678 16584
rect 8386 16532 8392 16584
rect 8444 16532 8450 16584
rect 9140 16572 9168 16612
rect 10060 16612 11060 16640
rect 10060 16572 10088 16612
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 9140 16544 10088 16572
rect 6730 16504 6736 16516
rect 6670 16476 6736 16504
rect 6730 16464 6736 16476
rect 6788 16464 6794 16516
rect 7282 16464 7288 16516
rect 7340 16464 7346 16516
rect 9300 16507 9358 16513
rect 9300 16473 9312 16507
rect 9346 16504 9358 16507
rect 9766 16504 9772 16516
rect 9346 16476 9772 16504
rect 9346 16473 9358 16476
rect 9300 16467 9358 16473
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 3053 16439 3111 16445
rect 3053 16436 3065 16439
rect 2832 16408 3065 16436
rect 2832 16396 2838 16408
rect 3053 16405 3065 16408
rect 3099 16405 3111 16439
rect 3053 16399 3111 16405
rect 4249 16439 4307 16445
rect 4249 16405 4261 16439
rect 4295 16405 4307 16439
rect 4249 16399 4307 16405
rect 4709 16439 4767 16445
rect 4709 16405 4721 16439
rect 4755 16436 4767 16439
rect 5166 16436 5172 16448
rect 4755 16408 5172 16436
rect 4755 16405 4767 16408
rect 4709 16399 4767 16405
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 10413 16439 10471 16445
rect 10413 16436 10425 16439
rect 9456 16408 10425 16436
rect 9456 16396 9462 16408
rect 10413 16405 10425 16408
rect 10459 16405 10471 16439
rect 10413 16399 10471 16405
rect 1104 16346 16811 16368
rect 1104 16294 4836 16346
rect 4888 16294 4900 16346
rect 4952 16294 4964 16346
rect 5016 16294 5028 16346
rect 5080 16294 5092 16346
rect 5144 16294 8723 16346
rect 8775 16294 8787 16346
rect 8839 16294 8851 16346
rect 8903 16294 8915 16346
rect 8967 16294 8979 16346
rect 9031 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 16497 16346
rect 16549 16294 16561 16346
rect 16613 16294 16625 16346
rect 16677 16294 16689 16346
rect 16741 16294 16753 16346
rect 16805 16294 16811 16346
rect 1104 16272 16811 16294
rect 2130 16192 2136 16244
rect 2188 16192 2194 16244
rect 2593 16235 2651 16241
rect 2593 16201 2605 16235
rect 2639 16201 2651 16235
rect 2593 16195 2651 16201
rect 2317 16099 2375 16105
rect 2317 16065 2329 16099
rect 2363 16096 2375 16099
rect 2608 16096 2636 16195
rect 2682 16192 2688 16244
rect 2740 16232 2746 16244
rect 2740 16204 6408 16232
rect 2740 16192 2746 16204
rect 3053 16167 3111 16173
rect 3053 16133 3065 16167
rect 3099 16164 3111 16167
rect 3789 16167 3847 16173
rect 3789 16164 3801 16167
rect 3099 16136 3801 16164
rect 3099 16133 3111 16136
rect 3053 16127 3111 16133
rect 3789 16133 3801 16136
rect 3835 16133 3847 16167
rect 6270 16164 6276 16176
rect 5934 16136 6276 16164
rect 3789 16127 3847 16133
rect 6270 16124 6276 16136
rect 6328 16124 6334 16176
rect 2363 16068 2636 16096
rect 2363 16065 2375 16068
rect 2317 16059 2375 16065
rect 2774 16056 2780 16108
rect 2832 16096 2838 16108
rect 2961 16099 3019 16105
rect 2961 16096 2973 16099
rect 2832 16068 2973 16096
rect 2832 16056 2838 16068
rect 2961 16065 2973 16068
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 3694 16096 3700 16108
rect 3651 16068 3700 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 3694 16056 3700 16068
rect 3752 16056 3758 16108
rect 4433 16099 4491 16105
rect 4433 16096 4445 16099
rect 3804 16068 4445 16096
rect 3804 16040 3832 16068
rect 4433 16065 4445 16068
rect 4479 16065 4491 16099
rect 4433 16059 4491 16065
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 15997 3295 16031
rect 3237 15991 3295 15997
rect 3252 15960 3280 15991
rect 3418 15988 3424 16040
rect 3476 15988 3482 16040
rect 3786 15988 3792 16040
rect 3844 15988 3850 16040
rect 4154 15988 4160 16040
rect 4212 15988 4218 16040
rect 4706 15988 4712 16040
rect 4764 15988 4770 16040
rect 4172 15960 4200 15988
rect 3252 15932 4200 15960
rect 6178 15852 6184 15904
rect 6236 15852 6242 15904
rect 6380 15892 6408 16204
rect 6454 16192 6460 16244
rect 6512 16192 6518 16244
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 7009 16235 7067 16241
rect 7009 16232 7021 16235
rect 6788 16204 7021 16232
rect 6788 16192 6794 16204
rect 7009 16201 7021 16204
rect 7055 16201 7067 16235
rect 7009 16195 7067 16201
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 7469 16235 7527 16241
rect 7469 16232 7481 16235
rect 7340 16204 7481 16232
rect 7340 16192 7346 16204
rect 7469 16201 7481 16204
rect 7515 16201 7527 16235
rect 7469 16195 7527 16201
rect 8110 16192 8116 16244
rect 8168 16192 8174 16244
rect 8386 16192 8392 16244
rect 8444 16192 8450 16244
rect 9309 16235 9367 16241
rect 9309 16201 9321 16235
rect 9355 16232 9367 16235
rect 9398 16232 9404 16244
rect 9355 16204 9404 16232
rect 9355 16201 9367 16204
rect 9309 16195 9367 16201
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 9766 16192 9772 16244
rect 9824 16192 9830 16244
rect 11149 16235 11207 16241
rect 11149 16201 11161 16235
rect 11195 16201 11207 16235
rect 11149 16195 11207 16201
rect 13265 16235 13323 16241
rect 13265 16201 13277 16235
rect 13311 16232 13323 16235
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13311 16204 13737 16232
rect 13311 16201 13323 16204
rect 13265 16195 13323 16201
rect 13725 16201 13737 16204
rect 13771 16201 13783 16235
rect 13725 16195 13783 16201
rect 8128 16164 8156 16192
rect 11164 16164 11192 16195
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 6656 16136 8156 16164
rect 8312 16136 10456 16164
rect 11164 16136 11805 16164
rect 6656 16105 6684 16136
rect 6641 16099 6699 16105
rect 6641 16065 6653 16099
rect 6687 16065 6699 16099
rect 6641 16059 6699 16065
rect 6917 16099 6975 16105
rect 6917 16065 6929 16099
rect 6963 16065 6975 16099
rect 6917 16059 6975 16065
rect 6932 15960 6960 16059
rect 7650 16056 7656 16108
rect 7708 16056 7714 16108
rect 7926 16056 7932 16108
rect 7984 16096 7990 16108
rect 8312 16105 8340 16136
rect 10428 16108 10456 16136
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 11793 16127 11851 16133
rect 12250 16124 12256 16176
rect 12308 16124 12314 16176
rect 8297 16099 8355 16105
rect 8297 16096 8309 16099
rect 7984 16068 8309 16096
rect 7984 16056 7990 16068
rect 8297 16065 8309 16068
rect 8343 16065 8355 16099
rect 8297 16059 8355 16065
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 7944 15960 7972 16056
rect 9398 15988 9404 16040
rect 9456 15988 9462 16040
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 6932 15932 7972 15960
rect 8941 15963 8999 15969
rect 8941 15929 8953 15963
rect 8987 15960 8999 15963
rect 9968 15960 9996 16059
rect 10410 16056 10416 16108
rect 10468 16056 10474 16108
rect 11330 16056 11336 16108
rect 11388 16056 11394 16108
rect 11514 15988 11520 16040
rect 11572 15988 11578 16040
rect 13170 15988 13176 16040
rect 13228 16028 13234 16040
rect 13817 16031 13875 16037
rect 13817 16028 13829 16031
rect 13228 16000 13829 16028
rect 13228 15988 13234 16000
rect 13817 15997 13829 16000
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 8987 15932 9996 15960
rect 8987 15929 8999 15932
rect 8941 15923 8999 15929
rect 13722 15920 13728 15972
rect 13780 15960 13786 15972
rect 13924 15960 13952 15991
rect 13780 15932 13952 15960
rect 13780 15920 13786 15932
rect 8386 15892 8392 15904
rect 6380 15864 8392 15892
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 13354 15852 13360 15904
rect 13412 15852 13418 15904
rect 1104 15802 16652 15824
rect 1104 15750 2893 15802
rect 2945 15750 2957 15802
rect 3009 15750 3021 15802
rect 3073 15750 3085 15802
rect 3137 15750 3149 15802
rect 3201 15750 6780 15802
rect 6832 15750 6844 15802
rect 6896 15750 6908 15802
rect 6960 15750 6972 15802
rect 7024 15750 7036 15802
rect 7088 15750 10667 15802
rect 10719 15750 10731 15802
rect 10783 15750 10795 15802
rect 10847 15750 10859 15802
rect 10911 15750 10923 15802
rect 10975 15750 14554 15802
rect 14606 15750 14618 15802
rect 14670 15750 14682 15802
rect 14734 15750 14746 15802
rect 14798 15750 14810 15802
rect 14862 15750 16652 15802
rect 1104 15728 16652 15750
rect 3418 15648 3424 15700
rect 3476 15648 3482 15700
rect 4706 15648 4712 15700
rect 4764 15688 4770 15700
rect 5261 15691 5319 15697
rect 5261 15688 5273 15691
rect 4764 15660 5273 15688
rect 4764 15648 4770 15660
rect 5261 15657 5273 15660
rect 5307 15657 5319 15691
rect 5261 15651 5319 15657
rect 6270 15648 6276 15700
rect 6328 15648 6334 15700
rect 9398 15648 9404 15700
rect 9456 15648 9462 15700
rect 12250 15648 12256 15700
rect 12308 15648 12314 15700
rect 13354 15648 13360 15700
rect 13412 15648 13418 15700
rect 3436 15620 3464 15648
rect 3436 15592 5120 15620
rect 5092 15552 5120 15592
rect 5166 15580 5172 15632
rect 5224 15580 5230 15632
rect 10226 15620 10232 15632
rect 8956 15592 10232 15620
rect 8956 15552 8984 15592
rect 10226 15580 10232 15592
rect 10284 15620 10290 15632
rect 11882 15620 11888 15632
rect 10284 15592 11888 15620
rect 10284 15580 10290 15592
rect 11882 15580 11888 15592
rect 11940 15580 11946 15632
rect 5092 15524 8984 15552
rect 9033 15555 9091 15561
rect 9033 15521 9045 15555
rect 9079 15552 9091 15555
rect 9079 15524 9812 15552
rect 9079 15521 9091 15524
rect 9033 15515 9091 15521
rect 3694 15444 3700 15496
rect 3752 15444 3758 15496
rect 4890 15444 4896 15496
rect 4948 15444 4954 15496
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15453 5043 15487
rect 4985 15447 5043 15453
rect 3712 15416 3740 15444
rect 5000 15416 5028 15447
rect 5258 15444 5264 15496
rect 5316 15484 5322 15496
rect 5445 15487 5503 15493
rect 5445 15484 5457 15487
rect 5316 15456 5457 15484
rect 5316 15444 5322 15456
rect 5445 15453 5457 15456
rect 5491 15453 5503 15487
rect 5445 15447 5503 15453
rect 6181 15487 6239 15493
rect 6181 15453 6193 15487
rect 6227 15484 6239 15487
rect 7926 15484 7932 15496
rect 6227 15456 7932 15484
rect 6227 15453 6239 15456
rect 6181 15447 6239 15453
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 3712 15388 5028 15416
rect 9232 15360 9260 15447
rect 4890 15308 4896 15360
rect 4948 15348 4954 15360
rect 5442 15348 5448 15360
rect 4948 15320 5448 15348
rect 4948 15308 4954 15320
rect 5442 15308 5448 15320
rect 5500 15348 5506 15360
rect 8018 15348 8024 15360
rect 5500 15320 8024 15348
rect 5500 15308 5506 15320
rect 8018 15308 8024 15320
rect 8076 15308 8082 15360
rect 9214 15308 9220 15360
rect 9272 15308 9278 15360
rect 9784 15357 9812 15524
rect 12161 15487 12219 15493
rect 12161 15453 12173 15487
rect 12207 15453 12219 15487
rect 12161 15447 12219 15453
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15484 13047 15487
rect 13372 15484 13400 15648
rect 13035 15456 13400 15484
rect 14093 15487 14151 15493
rect 13035 15453 13047 15456
rect 12989 15447 13047 15453
rect 14093 15453 14105 15487
rect 14139 15484 14151 15487
rect 14366 15484 14372 15496
rect 14139 15456 14372 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 10410 15376 10416 15428
rect 10468 15416 10474 15428
rect 12176 15416 12204 15447
rect 14108 15416 14136 15447
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 10468 15388 14136 15416
rect 10468 15376 10474 15388
rect 9769 15351 9827 15357
rect 9769 15317 9781 15351
rect 9815 15348 9827 15351
rect 10042 15348 10048 15360
rect 9815 15320 10048 15348
rect 9815 15317 9827 15320
rect 9769 15311 9827 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 12805 15351 12863 15357
rect 12805 15317 12817 15351
rect 12851 15348 12863 15351
rect 13078 15348 13084 15360
rect 12851 15320 13084 15348
rect 12851 15317 12863 15320
rect 12805 15311 12863 15317
rect 13078 15308 13084 15320
rect 13136 15308 13142 15360
rect 14182 15308 14188 15360
rect 14240 15308 14246 15360
rect 1104 15258 16811 15280
rect 1104 15206 4836 15258
rect 4888 15206 4900 15258
rect 4952 15206 4964 15258
rect 5016 15206 5028 15258
rect 5080 15206 5092 15258
rect 5144 15206 8723 15258
rect 8775 15206 8787 15258
rect 8839 15206 8851 15258
rect 8903 15206 8915 15258
rect 8967 15206 8979 15258
rect 9031 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 16497 15258
rect 16549 15206 16561 15258
rect 16613 15206 16625 15258
rect 16677 15206 16689 15258
rect 16741 15206 16753 15258
rect 16805 15206 16811 15258
rect 1104 15184 16811 15206
rect 1486 15104 1492 15156
rect 1544 15144 1550 15156
rect 2314 15144 2320 15156
rect 1544 15116 2320 15144
rect 1544 15104 1550 15116
rect 2314 15104 2320 15116
rect 2372 15144 2378 15156
rect 2777 15147 2835 15153
rect 2777 15144 2789 15147
rect 2372 15116 2789 15144
rect 2372 15104 2378 15116
rect 2777 15113 2789 15116
rect 2823 15113 2835 15147
rect 2777 15107 2835 15113
rect 7377 15147 7435 15153
rect 7377 15113 7389 15147
rect 7423 15144 7435 15147
rect 7650 15144 7656 15156
rect 7423 15116 7656 15144
rect 7423 15113 7435 15116
rect 7377 15107 7435 15113
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 8294 15104 8300 15156
rect 8352 15104 8358 15156
rect 11333 15147 11391 15153
rect 9600 15116 11284 15144
rect 8312 15076 8340 15104
rect 9122 15076 9128 15088
rect 8036 15048 9128 15076
rect 1670 15017 1676 15020
rect 1664 14971 1676 15017
rect 1670 14968 1676 14971
rect 1728 14968 1734 15020
rect 7742 14968 7748 15020
rect 7800 14968 7806 15020
rect 1394 14900 1400 14952
rect 1452 14900 1458 14952
rect 8036 14949 8064 15048
rect 9122 15036 9128 15048
rect 9180 15036 9186 15088
rect 9306 15036 9312 15088
rect 9364 15076 9370 15088
rect 9600 15076 9628 15116
rect 9364 15048 9628 15076
rect 9364 15036 9370 15048
rect 9600 15017 9628 15048
rect 10502 15036 10508 15088
rect 10560 15036 10566 15088
rect 11256 15076 11284 15116
rect 11333 15113 11345 15147
rect 11379 15144 11391 15147
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11379 15116 11897 15144
rect 11379 15113 11391 15116
rect 11333 15107 11391 15113
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 11514 15076 11520 15088
rect 11256 15048 11520 15076
rect 11514 15036 11520 15048
rect 11572 15076 11578 15088
rect 12250 15076 12256 15088
rect 11572 15048 12256 15076
rect 11572 15036 11578 15048
rect 12250 15036 12256 15048
rect 12308 15076 12314 15088
rect 12308 15048 12434 15076
rect 12308 15036 12314 15048
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 15008 8355 15011
rect 9585 15011 9643 15017
rect 8343 14980 9536 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 7837 14943 7895 14949
rect 7837 14909 7849 14943
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 7852 14872 7880 14903
rect 8570 14872 8576 14884
rect 7852 14844 8576 14872
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 8389 14807 8447 14813
rect 8389 14804 8401 14807
rect 7524 14776 8401 14804
rect 7524 14764 7530 14776
rect 8389 14773 8401 14776
rect 8435 14773 8447 14807
rect 9508 14804 9536 14980
rect 9585 14977 9597 15011
rect 9631 14977 9643 15011
rect 12406 15008 12434 15048
rect 13078 15036 13084 15088
rect 13136 15076 13142 15088
rect 13173 15079 13231 15085
rect 13173 15076 13185 15079
rect 13136 15048 13185 15076
rect 13136 15036 13142 15048
rect 13173 15045 13185 15048
rect 13219 15045 13231 15079
rect 13173 15039 13231 15045
rect 14182 15036 14188 15088
rect 14240 15036 14246 15088
rect 12897 15011 12955 15017
rect 12897 15008 12909 15011
rect 9585 14971 9643 14977
rect 11256 14980 12112 15008
rect 12406 14980 12909 15008
rect 11256 14952 11284 14980
rect 9858 14900 9864 14952
rect 9916 14900 9922 14952
rect 11238 14900 11244 14952
rect 11296 14900 11302 14952
rect 11330 14900 11336 14952
rect 11388 14900 11394 14952
rect 11974 14900 11980 14952
rect 12032 14900 12038 14952
rect 12084 14949 12112 14980
rect 12897 14977 12909 14980
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 12069 14943 12127 14949
rect 12069 14909 12081 14943
rect 12115 14940 12127 14943
rect 13722 14940 13728 14952
rect 12115 14912 13728 14940
rect 12115 14909 12127 14912
rect 12069 14903 12127 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 11348 14872 11376 14900
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 11348 14844 11529 14872
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 13630 14804 13636 14816
rect 9508 14776 13636 14804
rect 8389 14767 8447 14773
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 14458 14764 14464 14816
rect 14516 14804 14522 14816
rect 14645 14807 14703 14813
rect 14645 14804 14657 14807
rect 14516 14776 14657 14804
rect 14516 14764 14522 14776
rect 14645 14773 14657 14776
rect 14691 14773 14703 14807
rect 14645 14767 14703 14773
rect 1104 14714 16652 14736
rect 1104 14662 2893 14714
rect 2945 14662 2957 14714
rect 3009 14662 3021 14714
rect 3073 14662 3085 14714
rect 3137 14662 3149 14714
rect 3201 14662 6780 14714
rect 6832 14662 6844 14714
rect 6896 14662 6908 14714
rect 6960 14662 6972 14714
rect 7024 14662 7036 14714
rect 7088 14662 10667 14714
rect 10719 14662 10731 14714
rect 10783 14662 10795 14714
rect 10847 14662 10859 14714
rect 10911 14662 10923 14714
rect 10975 14662 14554 14714
rect 14606 14662 14618 14714
rect 14670 14662 14682 14714
rect 14734 14662 14746 14714
rect 14798 14662 14810 14714
rect 14862 14662 16652 14714
rect 1104 14640 16652 14662
rect 1670 14560 1676 14612
rect 1728 14560 1734 14612
rect 7377 14603 7435 14609
rect 2608 14572 7328 14600
rect 1394 14424 1400 14476
rect 1452 14464 1458 14476
rect 2608 14473 2636 14572
rect 5166 14492 5172 14544
rect 5224 14492 5230 14544
rect 5261 14535 5319 14541
rect 5261 14501 5273 14535
rect 5307 14532 5319 14535
rect 7300 14532 7328 14572
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 7742 14600 7748 14612
rect 7423 14572 7748 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 9769 14603 9827 14609
rect 9769 14569 9781 14603
rect 9815 14600 9827 14603
rect 9858 14600 9864 14612
rect 9815 14572 9864 14600
rect 9815 14569 9827 14572
rect 9769 14563 9827 14569
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 10689 14603 10747 14609
rect 10689 14600 10701 14603
rect 10560 14572 10701 14600
rect 10560 14560 10566 14572
rect 10689 14569 10701 14572
rect 10735 14569 10747 14603
rect 10689 14563 10747 14569
rect 13170 14560 13176 14612
rect 13228 14560 13234 14612
rect 8294 14532 8300 14544
rect 5307 14504 5764 14532
rect 7300 14504 8300 14532
rect 5307 14501 5319 14504
rect 5261 14495 5319 14501
rect 2593 14467 2651 14473
rect 1452 14436 2544 14464
rect 1452 14424 1458 14436
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14396 1915 14399
rect 1903 14368 1992 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 1964 14269 1992 14368
rect 2314 14356 2320 14408
rect 2372 14356 2378 14408
rect 2516 14396 2544 14436
rect 2593 14433 2605 14467
rect 2639 14433 2651 14467
rect 3786 14464 3792 14476
rect 2593 14427 2651 14433
rect 3068 14436 3792 14464
rect 3068 14396 3096 14436
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 5736 14464 5764 14504
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 8941 14535 8999 14541
rect 8941 14501 8953 14535
rect 8987 14501 8999 14535
rect 8941 14495 8999 14501
rect 5905 14467 5963 14473
rect 5905 14464 5917 14467
rect 4816 14436 5580 14464
rect 5736 14436 5917 14464
rect 2516 14368 3096 14396
rect 3142 14356 3148 14408
rect 3200 14356 3206 14408
rect 3326 14356 3332 14408
rect 3384 14356 3390 14408
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 3694 14396 3700 14408
rect 3467 14368 3700 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 3694 14356 3700 14368
rect 3752 14356 3758 14408
rect 3804 14396 3832 14424
rect 4816 14396 4844 14436
rect 3804 14368 4844 14396
rect 4890 14356 4896 14408
rect 4948 14396 4954 14408
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 4948 14368 5457 14396
rect 4948 14356 4954 14368
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 5552 14396 5580 14436
rect 5905 14433 5917 14436
rect 5951 14433 5963 14467
rect 5905 14427 5963 14433
rect 5626 14396 5632 14408
rect 5552 14368 5632 14396
rect 5445 14359 5503 14365
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14396 7527 14399
rect 7650 14396 7656 14408
rect 7515 14368 7656 14396
rect 7515 14365 7527 14368
rect 7469 14359 7527 14365
rect 7650 14356 7656 14368
rect 7708 14396 7714 14408
rect 7926 14396 7932 14408
rect 7708 14368 7932 14396
rect 7708 14356 7714 14368
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14396 8079 14399
rect 8956 14396 8984 14495
rect 10410 14492 10416 14544
rect 10468 14492 10474 14544
rect 9582 14424 9588 14476
rect 9640 14424 9646 14476
rect 8067 14368 8984 14396
rect 8067 14365 8079 14368
rect 8021 14359 8079 14365
rect 9398 14356 9404 14408
rect 9456 14356 9462 14408
rect 9950 14356 9956 14408
rect 10008 14356 10014 14408
rect 10428 14396 10456 14492
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11793 14467 11851 14473
rect 11793 14464 11805 14467
rect 11112 14436 11805 14464
rect 11112 14424 11118 14436
rect 11793 14433 11805 14436
rect 11839 14433 11851 14467
rect 11793 14427 11851 14433
rect 13722 14424 13728 14476
rect 13780 14464 13786 14476
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 13780 14436 14657 14464
rect 13780 14424 13786 14436
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 10597 14399 10655 14405
rect 10597 14396 10609 14399
rect 10428 14368 10609 14396
rect 10597 14365 10609 14368
rect 10643 14365 10655 14399
rect 10597 14359 10655 14365
rect 14458 14356 14464 14408
rect 14516 14356 14522 14408
rect 4034 14331 4092 14337
rect 4034 14328 4046 14331
rect 2976 14300 4046 14328
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14229 2007 14263
rect 1949 14223 2007 14229
rect 2409 14263 2467 14269
rect 2409 14229 2421 14263
rect 2455 14260 2467 14263
rect 2590 14260 2596 14272
rect 2455 14232 2596 14260
rect 2455 14229 2467 14232
rect 2409 14223 2467 14229
rect 2590 14220 2596 14232
rect 2648 14220 2654 14272
rect 2976 14269 3004 14300
rect 4034 14297 4046 14300
rect 4080 14297 4092 14331
rect 7561 14331 7619 14337
rect 7561 14328 7573 14331
rect 7130 14300 7573 14328
rect 4034 14291 4092 14297
rect 7561 14297 7573 14300
rect 7607 14297 7619 14331
rect 7561 14291 7619 14297
rect 7668 14300 7972 14328
rect 2961 14263 3019 14269
rect 2961 14229 2973 14263
rect 3007 14229 3019 14263
rect 2961 14223 3019 14229
rect 3602 14220 3608 14272
rect 3660 14220 3666 14272
rect 3878 14220 3884 14272
rect 3936 14260 3942 14272
rect 7668 14260 7696 14300
rect 3936 14232 7696 14260
rect 3936 14220 3942 14232
rect 7834 14220 7840 14272
rect 7892 14220 7898 14272
rect 7944 14260 7972 14300
rect 8570 14288 8576 14340
rect 8628 14328 8634 14340
rect 9309 14331 9367 14337
rect 9309 14328 9321 14331
rect 8628 14300 9321 14328
rect 8628 14288 8634 14300
rect 9309 14297 9321 14300
rect 9355 14297 9367 14331
rect 11514 14328 11520 14340
rect 9309 14291 9367 14297
rect 9416 14300 11520 14328
rect 9416 14260 9444 14300
rect 11514 14288 11520 14300
rect 11572 14288 11578 14340
rect 12060 14331 12118 14337
rect 12060 14297 12072 14331
rect 12106 14328 12118 14331
rect 12342 14328 12348 14340
rect 12106 14300 12348 14328
rect 12106 14297 12118 14300
rect 12060 14291 12118 14297
rect 12342 14288 12348 14300
rect 12400 14288 12406 14340
rect 12452 14300 16252 14328
rect 7944 14232 9444 14260
rect 10502 14220 10508 14272
rect 10560 14260 10566 14272
rect 12452 14260 12480 14300
rect 16224 14272 16252 14300
rect 10560 14232 12480 14260
rect 10560 14220 10566 14232
rect 14090 14220 14096 14272
rect 14148 14220 14154 14272
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 14553 14263 14611 14269
rect 14553 14260 14565 14263
rect 14332 14232 14565 14260
rect 14332 14220 14338 14232
rect 14553 14229 14565 14232
rect 14599 14229 14611 14263
rect 14553 14223 14611 14229
rect 16206 14220 16212 14272
rect 16264 14220 16270 14272
rect 1104 14170 16811 14192
rect 1104 14118 4836 14170
rect 4888 14118 4900 14170
rect 4952 14118 4964 14170
rect 5016 14118 5028 14170
rect 5080 14118 5092 14170
rect 5144 14118 8723 14170
rect 8775 14118 8787 14170
rect 8839 14118 8851 14170
rect 8903 14118 8915 14170
rect 8967 14118 8979 14170
rect 9031 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 16497 14170
rect 16549 14118 16561 14170
rect 16613 14118 16625 14170
rect 16677 14118 16689 14170
rect 16741 14118 16753 14170
rect 16805 14118 16811 14170
rect 1104 14096 16811 14118
rect 1762 14016 1768 14068
rect 1820 14056 1826 14068
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 1820 14028 1869 14056
rect 1820 14016 1826 14028
rect 1857 14025 1869 14028
rect 1903 14025 1915 14059
rect 1857 14019 1915 14025
rect 2225 14059 2283 14065
rect 2225 14025 2237 14059
rect 2271 14025 2283 14059
rect 2225 14019 2283 14025
rect 2685 14059 2743 14065
rect 2685 14025 2697 14059
rect 2731 14056 2743 14059
rect 2774 14056 2780 14068
rect 2731 14028 2780 14056
rect 2731 14025 2743 14028
rect 2685 14019 2743 14025
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 2240 13920 2268 14019
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 3421 14059 3479 14065
rect 3421 14056 3433 14059
rect 3200 14028 3433 14056
rect 3200 14016 3206 14028
rect 3421 14025 3433 14028
rect 3467 14025 3479 14059
rect 3421 14019 3479 14025
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 3881 14059 3939 14065
rect 3881 14056 3893 14059
rect 3660 14028 3893 14056
rect 3660 14016 3666 14028
rect 3881 14025 3893 14028
rect 3927 14025 3939 14059
rect 3881 14019 3939 14025
rect 4341 14059 4399 14065
rect 4341 14025 4353 14059
rect 4387 14056 4399 14059
rect 4706 14056 4712 14068
rect 4387 14028 4712 14056
rect 4387 14025 4399 14028
rect 4341 14019 4399 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 5166 14056 5172 14068
rect 4847 14028 5172 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 3789 13991 3847 13997
rect 3789 13957 3801 13991
rect 3835 13988 3847 13991
rect 4816 13988 4844 14019
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 5721 14059 5779 14065
rect 5721 14025 5733 14059
rect 5767 14025 5779 14059
rect 5721 14019 5779 14025
rect 5736 13988 5764 14019
rect 7834 14016 7840 14068
rect 7892 14016 7898 14068
rect 8570 14016 8576 14068
rect 8628 14056 8634 14068
rect 8849 14059 8907 14065
rect 8849 14056 8861 14059
rect 8628 14028 8861 14056
rect 8628 14016 8634 14028
rect 8849 14025 8861 14028
rect 8895 14025 8907 14059
rect 8849 14019 8907 14025
rect 9309 14059 9367 14065
rect 9309 14025 9321 14059
rect 9355 14056 9367 14059
rect 9398 14056 9404 14068
rect 9355 14028 9404 14056
rect 9355 14025 9367 14028
rect 9309 14019 9367 14025
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9950 14016 9956 14068
rect 10008 14016 10014 14068
rect 12342 14016 12348 14068
rect 12400 14016 12406 14068
rect 13170 14016 13176 14068
rect 13228 14016 13234 14068
rect 14090 14016 14096 14068
rect 14148 14016 14154 14068
rect 14366 14016 14372 14068
rect 14424 14016 14430 14068
rect 16206 14016 16212 14068
rect 16264 14016 16270 14068
rect 3835 13960 4844 13988
rect 4908 13960 5764 13988
rect 7736 13991 7794 13997
rect 3835 13957 3847 13960
rect 3789 13951 3847 13957
rect 2087 13892 2268 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2590 13880 2596 13932
rect 2648 13920 2654 13932
rect 2648 13892 4200 13920
rect 2648 13880 2654 13892
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 2869 13815 2927 13821
rect 2884 13784 2912 13815
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 3878 13852 3884 13864
rect 3476 13824 3884 13852
rect 3476 13812 3482 13824
rect 3878 13812 3884 13824
rect 3936 13812 3942 13864
rect 4062 13812 4068 13864
rect 4120 13812 4126 13864
rect 4172 13852 4200 13892
rect 4706 13880 4712 13932
rect 4764 13880 4770 13932
rect 4908 13920 4936 13960
rect 7736 13957 7748 13991
rect 7782 13988 7794 13991
rect 7852 13988 7880 14016
rect 11422 13988 11428 14000
rect 7782 13960 7880 13988
rect 9048 13960 11428 13988
rect 7782 13957 7794 13960
rect 7736 13951 7794 13957
rect 4816 13892 4936 13920
rect 4816 13852 4844 13892
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 7466 13920 7472 13932
rect 5684 13892 7472 13920
rect 5684 13880 5690 13892
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 9048 13929 9076 13960
rect 11422 13948 11428 13960
rect 11480 13948 11486 14000
rect 12069 13991 12127 13997
rect 12069 13957 12081 13991
rect 12115 13988 12127 13991
rect 13188 13988 13216 14016
rect 12115 13960 13216 13988
rect 12115 13957 12127 13960
rect 12069 13951 12127 13957
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13889 9091 13923
rect 9033 13883 9091 13889
rect 9125 13923 9183 13929
rect 9125 13889 9137 13923
rect 9171 13920 9183 13923
rect 9171 13892 9260 13920
rect 9171 13889 9183 13892
rect 9125 13883 9183 13889
rect 9232 13864 9260 13892
rect 10318 13880 10324 13932
rect 10376 13880 10382 13932
rect 10413 13923 10471 13929
rect 10413 13889 10425 13923
rect 10459 13920 10471 13923
rect 11054 13920 11060 13932
rect 10459 13892 11060 13920
rect 10459 13889 10471 13892
rect 10413 13883 10471 13889
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 11514 13880 11520 13932
rect 11572 13920 11578 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11572 13892 11805 13920
rect 11572 13880 11578 13892
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 4172 13824 4844 13852
rect 4985 13855 5043 13861
rect 4985 13821 4997 13855
rect 5031 13821 5043 13855
rect 4985 13815 5043 13821
rect 5000 13784 5028 13815
rect 5258 13812 5264 13864
rect 5316 13812 5322 13864
rect 9214 13812 9220 13864
rect 9272 13812 9278 13864
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13821 10563 13855
rect 11992 13852 12020 13883
rect 12158 13880 12164 13932
rect 12216 13880 12222 13932
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13153 13923 13211 13929
rect 13153 13920 13165 13923
rect 13044 13892 13165 13920
rect 13044 13880 13050 13892
rect 13153 13889 13165 13892
rect 13199 13889 13211 13923
rect 13153 13883 13211 13889
rect 12066 13852 12072 13864
rect 11992 13824 12072 13852
rect 10505 13815 10563 13821
rect 2884 13756 5672 13784
rect 5644 13728 5672 13756
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 10520 13784 10548 13815
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 12250 13812 12256 13864
rect 12308 13852 12314 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12308 13824 12909 13852
rect 12308 13812 12314 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 14108 13852 14136 14016
rect 14384 13929 14412 14016
rect 14461 13991 14519 13997
rect 14461 13957 14473 13991
rect 14507 13988 14519 13991
rect 15378 13988 15384 14000
rect 14507 13960 15384 13988
rect 14507 13957 14519 13960
rect 14461 13951 14519 13957
rect 15378 13948 15384 13960
rect 15436 13948 15442 14000
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16071 13892 16620 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 14844 13852 14872 13883
rect 16592 13864 16620 13892
rect 14108 13824 14872 13852
rect 12897 13815 12955 13821
rect 11238 13784 11244 13796
rect 9180 13756 11244 13784
rect 9180 13744 9186 13756
rect 11238 13744 11244 13756
rect 11296 13744 11302 13796
rect 5626 13676 5632 13728
rect 5684 13676 5690 13728
rect 12912 13716 12940 13815
rect 16574 13812 16580 13864
rect 16632 13812 16638 13864
rect 14366 13744 14372 13796
rect 14424 13784 14430 13796
rect 14645 13787 14703 13793
rect 14645 13784 14657 13787
rect 14424 13756 14657 13784
rect 14424 13744 14430 13756
rect 14645 13753 14657 13756
rect 14691 13753 14703 13787
rect 14645 13747 14703 13753
rect 13814 13716 13820 13728
rect 12912 13688 13820 13716
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14274 13676 14280 13728
rect 14332 13676 14338 13728
rect 1104 13626 16652 13648
rect 1104 13574 2893 13626
rect 2945 13574 2957 13626
rect 3009 13574 3021 13626
rect 3073 13574 3085 13626
rect 3137 13574 3149 13626
rect 3201 13574 6780 13626
rect 6832 13574 6844 13626
rect 6896 13574 6908 13626
rect 6960 13574 6972 13626
rect 7024 13574 7036 13626
rect 7088 13574 10667 13626
rect 10719 13574 10731 13626
rect 10783 13574 10795 13626
rect 10847 13574 10859 13626
rect 10911 13574 10923 13626
rect 10975 13574 14554 13626
rect 14606 13574 14618 13626
rect 14670 13574 14682 13626
rect 14734 13574 14746 13626
rect 14798 13574 14810 13626
rect 14862 13574 16652 13626
rect 1104 13552 16652 13574
rect 5077 13515 5135 13521
rect 5077 13481 5089 13515
rect 5123 13512 5135 13515
rect 5258 13512 5264 13524
rect 5123 13484 5264 13512
rect 5123 13481 5135 13484
rect 5077 13475 5135 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 10318 13472 10324 13524
rect 10376 13512 10382 13524
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10376 13484 10701 13512
rect 10376 13472 10382 13484
rect 10689 13481 10701 13484
rect 10735 13481 10747 13515
rect 10689 13475 10747 13481
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 12161 13515 12219 13521
rect 12161 13512 12173 13515
rect 11112 13484 12173 13512
rect 11112 13472 11118 13484
rect 12161 13481 12173 13484
rect 12207 13481 12219 13515
rect 12161 13475 12219 13481
rect 12897 13515 12955 13521
rect 12897 13481 12909 13515
rect 12943 13512 12955 13515
rect 12986 13512 12992 13524
rect 12943 13484 12992 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 3344 13416 5672 13444
rect 3344 13385 3372 13416
rect 5644 13388 5672 13416
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13345 3387 13379
rect 3329 13339 3387 13345
rect 4706 13336 4712 13388
rect 4764 13336 4770 13388
rect 5626 13336 5632 13388
rect 5684 13336 5690 13388
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13376 8999 13379
rect 9306 13376 9312 13388
rect 8987 13348 9312 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 13814 13336 13820 13388
rect 13872 13376 13878 13388
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 13872 13348 14105 13376
rect 13872 13336 13878 13348
rect 14093 13345 14105 13348
rect 14139 13345 14151 13379
rect 14093 13339 14151 13345
rect 14366 13336 14372 13388
rect 14424 13336 14430 13388
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 6178 13308 6184 13320
rect 4847 13280 6184 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 7282 13268 7288 13320
rect 7340 13308 7346 13320
rect 8113 13311 8171 13317
rect 8113 13308 8125 13311
rect 7340 13280 8125 13308
rect 7340 13268 7346 13280
rect 8113 13277 8125 13280
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13277 10839 13311
rect 10781 13271 10839 13277
rect 9217 13243 9275 13249
rect 9217 13240 9229 13243
rect 7944 13212 9229 13240
rect 2682 13132 2688 13184
rect 2740 13132 2746 13184
rect 3050 13132 3056 13184
rect 3108 13132 3114 13184
rect 3145 13175 3203 13181
rect 3145 13141 3157 13175
rect 3191 13172 3203 13175
rect 3326 13172 3332 13184
rect 3191 13144 3332 13172
rect 3191 13141 3203 13144
rect 3145 13135 3203 13141
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 7944 13181 7972 13212
rect 9217 13209 9229 13212
rect 9263 13209 9275 13243
rect 9217 13203 9275 13209
rect 9490 13200 9496 13252
rect 9548 13240 9554 13252
rect 9548 13212 9706 13240
rect 9548 13200 9554 13212
rect 7929 13175 7987 13181
rect 7929 13141 7941 13175
rect 7975 13141 7987 13175
rect 7929 13135 7987 13141
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 10796 13172 10824 13271
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 11480 13280 12357 13308
rect 11480 13268 11486 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 12345 13271 12403 13277
rect 12452 13280 12725 13308
rect 11048 13243 11106 13249
rect 11048 13209 11060 13243
rect 11094 13240 11106 13243
rect 11330 13240 11336 13252
rect 11094 13212 11336 13240
rect 11094 13209 11106 13212
rect 11048 13203 11106 13209
rect 11330 13200 11336 13212
rect 11388 13200 11394 13252
rect 11882 13200 11888 13252
rect 11940 13240 11946 13252
rect 12158 13240 12164 13252
rect 11940 13212 12164 13240
rect 11940 13200 11946 13212
rect 12158 13200 12164 13212
rect 12216 13240 12222 13252
rect 12452 13240 12480 13280
rect 12713 13277 12725 13280
rect 12759 13277 12771 13311
rect 12713 13271 12771 13277
rect 12216 13212 12480 13240
rect 12529 13243 12587 13249
rect 12216 13200 12222 13212
rect 12529 13209 12541 13243
rect 12575 13209 12587 13243
rect 12529 13203 12587 13209
rect 12621 13243 12679 13249
rect 12621 13209 12633 13243
rect 12667 13240 12679 13243
rect 14274 13240 14280 13252
rect 12667 13212 14280 13240
rect 12667 13209 12679 13212
rect 12621 13203 12679 13209
rect 11146 13172 11152 13184
rect 10008 13144 11152 13172
rect 10008 13132 10014 13144
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12544 13172 12572 13203
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 15378 13200 15384 13252
rect 15436 13200 15442 13252
rect 12492 13144 12572 13172
rect 12492 13132 12498 13144
rect 15838 13132 15844 13184
rect 15896 13132 15902 13184
rect 1104 13082 16811 13104
rect 1104 13030 4836 13082
rect 4888 13030 4900 13082
rect 4952 13030 4964 13082
rect 5016 13030 5028 13082
rect 5080 13030 5092 13082
rect 5144 13030 8723 13082
rect 8775 13030 8787 13082
rect 8839 13030 8851 13082
rect 8903 13030 8915 13082
rect 8967 13030 8979 13082
rect 9031 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 16497 13082
rect 16549 13030 16561 13082
rect 16613 13030 16625 13082
rect 16677 13030 16689 13082
rect 16741 13030 16753 13082
rect 16805 13030 16811 13082
rect 1104 13008 16811 13030
rect 2593 12971 2651 12977
rect 2593 12937 2605 12971
rect 2639 12937 2651 12971
rect 2593 12931 2651 12937
rect 4617 12971 4675 12977
rect 4617 12937 4629 12971
rect 4663 12968 4675 12971
rect 4706 12968 4712 12980
rect 4663 12940 4712 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 2608 12900 2636 12931
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 6178 12968 6184 12980
rect 5859 12940 6184 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8352 12940 8769 12968
rect 8352 12928 8358 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 8757 12931 8815 12937
rect 9033 12971 9091 12977
rect 9033 12937 9045 12971
rect 9079 12968 9091 12971
rect 9122 12968 9128 12980
rect 9079 12940 9128 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 3145 12903 3203 12909
rect 3145 12900 3157 12903
rect 2608 12872 3157 12900
rect 3145 12869 3157 12872
rect 3191 12869 3203 12903
rect 3145 12863 3203 12869
rect 4154 12860 4160 12912
rect 4212 12860 4218 12912
rect 7098 12860 7104 12912
rect 7156 12860 7162 12912
rect 8570 12860 8576 12912
rect 8628 12860 8634 12912
rect 1489 12835 1547 12841
rect 1489 12801 1501 12835
rect 1535 12801 1547 12835
rect 1489 12795 1547 12801
rect 1504 12764 1532 12795
rect 2314 12792 2320 12844
rect 2372 12792 2378 12844
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2740 12804 2789 12832
rect 2740 12792 2746 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 2866 12792 2872 12844
rect 2924 12792 2930 12844
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 3510 12764 3516 12776
rect 1504 12736 3516 12764
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 5902 12724 5908 12776
rect 5960 12724 5966 12776
rect 6089 12767 6147 12773
rect 6089 12733 6101 12767
rect 6135 12764 6147 12767
rect 6135 12736 6316 12764
rect 6135 12733 6147 12736
rect 6089 12727 6147 12733
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 2455 12668 2820 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 2792 12640 2820 12668
rect 1578 12588 1584 12640
rect 1636 12588 1642 12640
rect 2774 12588 2780 12640
rect 2832 12588 2838 12640
rect 5445 12631 5503 12637
rect 5445 12597 5457 12631
rect 5491 12628 5503 12631
rect 5718 12628 5724 12640
rect 5491 12600 5724 12628
rect 5491 12597 5503 12600
rect 5445 12591 5503 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 6288 12628 6316 12736
rect 6362 12724 6368 12776
rect 6420 12724 6426 12776
rect 6638 12724 6644 12776
rect 6696 12724 6702 12776
rect 7926 12764 7932 12776
rect 7668 12736 7932 12764
rect 7668 12628 7696 12736
rect 7926 12724 7932 12736
rect 7984 12764 7990 12776
rect 9048 12764 9076 12931
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9490 12928 9496 12980
rect 9548 12928 9554 12980
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 10284 12940 10824 12968
rect 10284 12928 10290 12940
rect 10410 12900 10416 12912
rect 9416 12872 10416 12900
rect 9416 12841 9444 12872
rect 10410 12860 10416 12872
rect 10468 12900 10474 12912
rect 10505 12903 10563 12909
rect 10505 12900 10517 12903
rect 10468 12872 10517 12900
rect 10468 12860 10474 12872
rect 10505 12869 10517 12872
rect 10551 12869 10563 12903
rect 10505 12863 10563 12869
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 10226 12792 10232 12844
rect 10284 12792 10290 12844
rect 10796 12841 10824 12940
rect 10980 12940 11192 12968
rect 10980 12909 11008 12940
rect 10965 12903 11023 12909
rect 10965 12869 10977 12903
rect 11011 12869 11023 12903
rect 10965 12863 11023 12869
rect 11054 12860 11060 12912
rect 11112 12860 11118 12912
rect 11164 12900 11192 12940
rect 11330 12928 11336 12980
rect 11388 12928 11394 12980
rect 12434 12968 12440 12980
rect 12176 12940 12440 12968
rect 11790 12900 11796 12912
rect 11164 12872 11796 12900
rect 11790 12860 11796 12872
rect 11848 12900 11854 12912
rect 12066 12900 12072 12912
rect 11848 12872 12072 12900
rect 11848 12860 11854 12872
rect 12066 12860 12072 12872
rect 12124 12900 12130 12912
rect 12176 12909 12204 12940
rect 12434 12928 12440 12940
rect 12492 12928 12498 12980
rect 13265 12971 13323 12977
rect 13265 12937 13277 12971
rect 13311 12968 13323 12971
rect 15838 12968 15844 12980
rect 13311 12940 15844 12968
rect 13311 12937 13323 12940
rect 13265 12931 13323 12937
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 12124 12872 12173 12900
rect 12124 12860 12130 12872
rect 12161 12869 12173 12872
rect 12207 12869 12219 12903
rect 12161 12863 12219 12869
rect 12253 12903 12311 12909
rect 12253 12869 12265 12903
rect 12299 12900 12311 12903
rect 13354 12900 13360 12912
rect 12299 12872 13360 12900
rect 12299 12869 12311 12872
rect 12253 12863 12311 12869
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 13722 12900 13728 12912
rect 13556 12872 13728 12900
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11882 12832 11888 12844
rect 11195 12804 11888 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 12345 12835 12403 12841
rect 12345 12801 12357 12835
rect 12391 12801 12403 12835
rect 12345 12795 12403 12801
rect 7984 12736 9076 12764
rect 7984 12724 7990 12736
rect 8205 12699 8263 12705
rect 8205 12665 8217 12699
rect 8251 12696 8263 12699
rect 8662 12696 8668 12708
rect 8251 12668 8668 12696
rect 8251 12665 8263 12668
rect 8205 12659 8263 12665
rect 8662 12656 8668 12668
rect 8720 12656 8726 12708
rect 6288 12600 7696 12628
rect 8110 12588 8116 12640
rect 8168 12588 8174 12640
rect 8386 12588 8392 12640
rect 8444 12628 8450 12640
rect 8573 12631 8631 12637
rect 8573 12628 8585 12631
rect 8444 12600 8585 12628
rect 8444 12588 8450 12600
rect 8573 12597 8585 12600
rect 8619 12597 8631 12631
rect 8573 12591 8631 12597
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 11992 12628 12020 12795
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12360 12764 12388 12795
rect 13556 12773 13584 12872
rect 13722 12860 13728 12872
rect 13780 12860 13786 12912
rect 13814 12860 13820 12912
rect 13872 12900 13878 12912
rect 13872 12872 14044 12900
rect 13872 12860 13878 12872
rect 13630 12792 13636 12844
rect 13688 12792 13694 12844
rect 14016 12841 14044 12872
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 12216 12736 12388 12764
rect 13541 12767 13599 12773
rect 12216 12724 12222 12736
rect 13541 12733 13553 12767
rect 13587 12733 13599 12767
rect 13648 12764 13676 12792
rect 13725 12767 13783 12773
rect 13725 12764 13737 12767
rect 13648 12736 13737 12764
rect 13541 12727 13599 12733
rect 13725 12733 13737 12736
rect 13771 12764 13783 12767
rect 13906 12764 13912 12776
rect 13771 12736 13912 12764
rect 13771 12733 13783 12736
rect 13725 12727 13783 12733
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 10100 12600 12020 12628
rect 10100 12588 10106 12600
rect 12526 12588 12532 12640
rect 12584 12588 12590 12640
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13814 12628 13820 12640
rect 12943 12600 13820 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 1104 12538 16652 12560
rect 1104 12486 2893 12538
rect 2945 12486 2957 12538
rect 3009 12486 3021 12538
rect 3073 12486 3085 12538
rect 3137 12486 3149 12538
rect 3201 12486 6780 12538
rect 6832 12486 6844 12538
rect 6896 12486 6908 12538
rect 6960 12486 6972 12538
rect 7024 12486 7036 12538
rect 7088 12486 10667 12538
rect 10719 12486 10731 12538
rect 10783 12486 10795 12538
rect 10847 12486 10859 12538
rect 10911 12486 10923 12538
rect 10975 12486 14554 12538
rect 14606 12486 14618 12538
rect 14670 12486 14682 12538
rect 14734 12486 14746 12538
rect 14798 12486 14810 12538
rect 14862 12486 16652 12538
rect 1104 12464 16652 12486
rect 2038 12424 2044 12436
rect 1504 12396 2044 12424
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1504 12288 1532 12396
rect 2038 12384 2044 12396
rect 2096 12424 2102 12436
rect 3145 12427 3203 12433
rect 2096 12396 2728 12424
rect 2096 12384 2102 12396
rect 2700 12368 2728 12396
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 3234 12424 3240 12436
rect 3191 12396 3240 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 4154 12424 4160 12436
rect 4019 12396 4160 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 5169 12427 5227 12433
rect 5169 12393 5181 12427
rect 5215 12424 5227 12427
rect 5350 12424 5356 12436
rect 5215 12396 5356 12424
rect 5215 12393 5227 12396
rect 5169 12387 5227 12393
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 5721 12427 5779 12433
rect 5721 12393 5733 12427
rect 5767 12424 5779 12427
rect 6638 12424 6644 12436
rect 5767 12396 6644 12424
rect 5767 12393 5779 12396
rect 5721 12387 5779 12393
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 6917 12427 6975 12433
rect 6917 12393 6929 12427
rect 6963 12424 6975 12427
rect 7098 12424 7104 12436
rect 6963 12396 7104 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7282 12384 7288 12436
rect 7340 12384 7346 12436
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 8536 12396 11836 12424
rect 8536 12384 8542 12396
rect 2682 12316 2688 12368
rect 2740 12316 2746 12368
rect 1443 12260 1532 12288
rect 1673 12291 1731 12297
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1673 12257 1685 12291
rect 1719 12288 1731 12291
rect 1762 12288 1768 12300
rect 1719 12260 1768 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 1762 12248 1768 12260
rect 1820 12248 1826 12300
rect 2314 12248 2320 12300
rect 2372 12288 2378 12300
rect 4893 12291 4951 12297
rect 2372 12260 3924 12288
rect 2372 12248 2378 12260
rect 3896 12232 3924 12260
rect 4893 12257 4905 12291
rect 4939 12288 4951 12291
rect 5534 12288 5540 12300
rect 4939 12260 5540 12288
rect 4939 12257 4951 12260
rect 4893 12251 4951 12257
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 7926 12248 7932 12300
rect 7984 12248 7990 12300
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12257 9275 12291
rect 11808 12288 11836 12396
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12161 12427 12219 12433
rect 12161 12424 12173 12427
rect 12032 12396 12173 12424
rect 12032 12384 12038 12396
rect 12161 12393 12173 12396
rect 12207 12393 12219 12427
rect 12161 12387 12219 12393
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 13412 12396 13645 12424
rect 13412 12384 13418 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 11808 12260 12388 12288
rect 9217 12251 9275 12257
rect 2774 12180 2780 12232
rect 2832 12180 2838 12232
rect 3878 12180 3884 12232
rect 3936 12180 3942 12232
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 4816 12084 4844 12183
rect 5902 12180 5908 12232
rect 5960 12180 5966 12232
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 7650 12220 7656 12232
rect 6871 12192 7656 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 9232 12220 9260 12251
rect 9766 12220 9772 12232
rect 9232 12192 9772 12220
rect 9766 12180 9772 12192
rect 9824 12220 9830 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 9824 12192 10793 12220
rect 9824 12180 9830 12192
rect 10781 12189 10793 12192
rect 10827 12220 10839 12223
rect 12250 12220 12256 12232
rect 10827 12192 12256 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 12360 12220 12388 12260
rect 12526 12229 12532 12232
rect 12360 12192 12434 12220
rect 8110 12152 8116 12164
rect 7668 12124 8116 12152
rect 7668 12093 7696 12124
rect 8110 12112 8116 12124
rect 8168 12112 8174 12164
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 9462 12155 9520 12161
rect 9462 12152 9474 12155
rect 9364 12124 9474 12152
rect 9364 12112 9370 12124
rect 9462 12121 9474 12124
rect 9508 12121 9520 12155
rect 9462 12115 9520 12121
rect 11048 12155 11106 12161
rect 11048 12121 11060 12155
rect 11094 12152 11106 12155
rect 12066 12152 12072 12164
rect 11094 12124 12072 12152
rect 11094 12121 11106 12124
rect 11048 12115 11106 12121
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 12406 12152 12434 12192
rect 12520 12183 12532 12229
rect 12526 12180 12532 12183
rect 12584 12180 12590 12232
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13872 12192 14289 12220
rect 13872 12180 13878 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 15746 12152 15752 12164
rect 12406 12124 15752 12152
rect 15746 12112 15752 12124
rect 15804 12112 15810 12164
rect 7653 12087 7711 12093
rect 7653 12084 7665 12087
rect 4816 12056 7665 12084
rect 7653 12053 7665 12056
rect 7699 12053 7711 12087
rect 7653 12047 7711 12053
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12084 7803 12087
rect 7926 12084 7932 12096
rect 7791 12056 7932 12084
rect 7791 12053 7803 12056
rect 7745 12047 7803 12053
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 10226 12044 10232 12096
rect 10284 12084 10290 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 10284 12056 10609 12084
rect 10284 12044 10290 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 14090 12044 14096 12096
rect 14148 12044 14154 12096
rect 1104 11994 16811 12016
rect 1104 11942 4836 11994
rect 4888 11942 4900 11994
rect 4952 11942 4964 11994
rect 5016 11942 5028 11994
rect 5080 11942 5092 11994
rect 5144 11942 8723 11994
rect 8775 11942 8787 11994
rect 8839 11942 8851 11994
rect 8903 11942 8915 11994
rect 8967 11942 8979 11994
rect 9031 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 16497 11994
rect 16549 11942 16561 11994
rect 16613 11942 16625 11994
rect 16677 11942 16689 11994
rect 16741 11942 16753 11994
rect 16805 11942 16811 11994
rect 1104 11920 16811 11942
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 9217 11883 9275 11889
rect 4028 11852 8064 11880
rect 4028 11840 4034 11852
rect 8036 11824 8064 11852
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 9306 11880 9312 11892
rect 9263 11852 9312 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 12066 11840 12072 11892
rect 12124 11840 12130 11892
rect 14090 11840 14096 11892
rect 14148 11840 14154 11892
rect 1872 11784 7604 11812
rect 1872 11552 1900 11784
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11744 2651 11747
rect 2774 11744 2780 11756
rect 2639 11716 2780 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6420 11716 6561 11744
rect 6420 11704 6426 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 6805 11747 6863 11753
rect 6805 11744 6817 11747
rect 6696 11716 6817 11744
rect 6696 11704 6702 11716
rect 6805 11713 6817 11716
rect 6851 11713 6863 11747
rect 6805 11707 6863 11713
rect 7576 11676 7604 11784
rect 8018 11772 8024 11824
rect 8076 11812 8082 11824
rect 8076 11784 11376 11812
rect 8076 11772 8082 11784
rect 11348 11756 11376 11784
rect 11698 11772 11704 11824
rect 11756 11772 11762 11824
rect 11793 11815 11851 11821
rect 11793 11781 11805 11815
rect 11839 11812 11851 11815
rect 11974 11812 11980 11824
rect 11839 11784 11980 11812
rect 11839 11781 11851 11784
rect 11793 11775 11851 11781
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 14001 11815 14059 11821
rect 14001 11781 14013 11815
rect 14047 11812 14059 11815
rect 14108 11812 14136 11840
rect 14047 11784 14136 11812
rect 14047 11781 14059 11784
rect 14001 11775 14059 11781
rect 15010 11772 15016 11824
rect 15068 11772 15074 11824
rect 9398 11704 9404 11756
rect 9456 11704 9462 11756
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11388 11716 11529 11744
rect 11388 11704 11394 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11882 11704 11888 11756
rect 11940 11704 11946 11756
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 13725 11747 13783 11753
rect 13725 11744 13737 11747
rect 12308 11716 13737 11744
rect 12308 11704 12314 11716
rect 13725 11713 13737 11716
rect 13771 11713 13783 11747
rect 13725 11707 13783 11713
rect 15838 11676 15844 11688
rect 7576 11648 15844 11676
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 9766 11608 9772 11620
rect 7852 11580 9772 11608
rect 1854 11500 1860 11552
rect 1912 11500 1918 11552
rect 2222 11500 2228 11552
rect 2280 11540 2286 11552
rect 2409 11543 2467 11549
rect 2409 11540 2421 11543
rect 2280 11512 2421 11540
rect 2280 11500 2286 11512
rect 2409 11509 2421 11512
rect 2455 11509 2467 11543
rect 2409 11503 2467 11509
rect 3878 11500 3884 11552
rect 3936 11540 3942 11552
rect 7852 11540 7880 11580
rect 9766 11568 9772 11580
rect 9824 11608 9830 11620
rect 10226 11608 10232 11620
rect 9824 11580 10232 11608
rect 9824 11568 9830 11580
rect 10226 11568 10232 11580
rect 10284 11568 10290 11620
rect 3936 11512 7880 11540
rect 3936 11500 3942 11512
rect 7926 11500 7932 11552
rect 7984 11500 7990 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 9582 11540 9588 11552
rect 8352 11512 9588 11540
rect 8352 11500 8358 11512
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 15470 11500 15476 11552
rect 15528 11500 15534 11552
rect 1104 11450 16652 11472
rect 1104 11398 2893 11450
rect 2945 11398 2957 11450
rect 3009 11398 3021 11450
rect 3073 11398 3085 11450
rect 3137 11398 3149 11450
rect 3201 11398 6780 11450
rect 6832 11398 6844 11450
rect 6896 11398 6908 11450
rect 6960 11398 6972 11450
rect 7024 11398 7036 11450
rect 7088 11398 10667 11450
rect 10719 11398 10731 11450
rect 10783 11398 10795 11450
rect 10847 11398 10859 11450
rect 10911 11398 10923 11450
rect 10975 11398 14554 11450
rect 14606 11398 14618 11450
rect 14670 11398 14682 11450
rect 14734 11398 14746 11450
rect 14798 11398 14810 11450
rect 14862 11398 16652 11450
rect 1104 11376 16652 11398
rect 3326 11296 3332 11348
rect 3384 11296 3390 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4120 11308 5672 11336
rect 4120 11296 4126 11308
rect 3970 11228 3976 11280
rect 4028 11228 4034 11280
rect 3786 11160 3792 11212
rect 3844 11200 3850 11212
rect 3988 11200 4016 11228
rect 3844 11172 4016 11200
rect 5644 11200 5672 11308
rect 5994 11296 6000 11348
rect 6052 11296 6058 11348
rect 8202 11296 8208 11348
rect 8260 11296 8266 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 8662 11336 8668 11348
rect 8619 11308 8668 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 8662 11296 8668 11308
rect 8720 11336 8726 11348
rect 9030 11336 9036 11348
rect 8720 11308 9036 11336
rect 8720 11296 8726 11308
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 9125 11339 9183 11345
rect 9125 11305 9137 11339
rect 9171 11336 9183 11339
rect 9398 11336 9404 11348
rect 9171 11308 9404 11336
rect 9171 11305 9183 11308
rect 9125 11299 9183 11305
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 14274 11336 14280 11348
rect 10980 11308 14280 11336
rect 6086 11228 6092 11280
rect 6144 11228 6150 11280
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 5644 11172 6745 11200
rect 3844 11160 3850 11172
rect 6733 11169 6745 11172
rect 6779 11200 6791 11203
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 6779 11172 7665 11200
rect 6779 11169 6791 11172
rect 6733 11163 6791 11169
rect 7653 11169 7665 11172
rect 7699 11200 7711 11203
rect 8220 11200 8248 11296
rect 8294 11228 8300 11280
rect 8352 11268 8358 11280
rect 8757 11271 8815 11277
rect 8757 11268 8769 11271
rect 8352 11240 8769 11268
rect 8352 11228 8358 11240
rect 8757 11237 8769 11240
rect 8803 11268 8815 11271
rect 9214 11268 9220 11280
rect 8803 11240 9220 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 8478 11200 8484 11212
rect 7699 11172 8248 11200
rect 8404 11172 8484 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 1854 11092 1860 11144
rect 1912 11092 1918 11144
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11132 2007 11135
rect 2038 11132 2044 11144
rect 1995 11104 2044 11132
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 2038 11092 2044 11104
rect 2096 11092 2102 11144
rect 2222 11141 2228 11144
rect 2216 11132 2228 11141
rect 2183 11104 2228 11132
rect 2216 11095 2228 11104
rect 2222 11092 2228 11095
rect 2280 11092 2286 11144
rect 3694 11092 3700 11144
rect 3752 11092 3758 11144
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 3712 11064 3740 11092
rect 3988 11064 4016 11095
rect 3712 11036 4016 11064
rect 1670 10956 1676 11008
rect 1728 10956 1734 11008
rect 4154 10956 4160 11008
rect 4212 10956 4218 11008
rect 4632 10996 4660 11095
rect 5994 11092 6000 11144
rect 6052 11132 6058 11144
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 6052 11104 6469 11132
rect 6052 11092 6058 11104
rect 6457 11101 6469 11104
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11132 7435 11135
rect 7926 11132 7932 11144
rect 7423 11104 7932 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 4706 11024 4712 11076
rect 4764 11064 4770 11076
rect 4862 11067 4920 11073
rect 4862 11064 4874 11067
rect 4764 11036 4874 11064
rect 4764 11024 4770 11036
rect 4862 11033 4874 11036
rect 4908 11033 4920 11067
rect 4862 11027 4920 11033
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 8404 11073 8432 11172
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 10980 11209 11008 11308
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 15470 11296 15476 11348
rect 15528 11296 15534 11348
rect 15838 11296 15844 11348
rect 15896 11296 15902 11348
rect 12161 11271 12219 11277
rect 12161 11237 12173 11271
rect 12207 11237 12219 11271
rect 12161 11231 12219 11237
rect 13633 11271 13691 11277
rect 13633 11237 13645 11271
rect 13679 11237 13691 11271
rect 13633 11231 13691 11237
rect 14369 11271 14427 11277
rect 14369 11237 14381 11271
rect 14415 11268 14427 11271
rect 15194 11268 15200 11280
rect 14415 11240 15200 11268
rect 14415 11237 14427 11240
rect 14369 11231 14427 11237
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 8628 11172 9689 11200
rect 8628 11160 8634 11172
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 10965 11203 11023 11209
rect 9677 11163 9735 11169
rect 9784 11172 10732 11200
rect 9784 11144 9812 11172
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9766 11132 9772 11144
rect 9539 11104 9772 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10502 11132 10508 11144
rect 9916 11104 10508 11132
rect 9916 11092 9922 11104
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 10704 11141 10732 11172
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11882 11160 11888 11212
rect 11940 11160 11946 11212
rect 12176 11200 12204 11231
rect 13648 11200 13676 11231
rect 15194 11228 15200 11240
rect 15252 11228 15258 11280
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 12176 11172 12388 11200
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11101 10747 11135
rect 10689 11095 10747 11101
rect 11609 11135 11667 11141
rect 11609 11101 11621 11135
rect 11655 11101 11667 11135
rect 11609 11095 11667 11101
rect 6549 11067 6607 11073
rect 6549 11064 6561 11067
rect 5868 11036 6561 11064
rect 5868 11024 5874 11036
rect 6549 11033 6561 11036
rect 6595 11033 6607 11067
rect 6549 11027 6607 11033
rect 8389 11067 8447 11073
rect 8389 11033 8401 11067
rect 8435 11064 8447 11067
rect 9398 11064 9404 11076
rect 8435 11036 9404 11064
rect 8435 11033 8447 11036
rect 8389 11027 8447 11033
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 9585 11067 9643 11073
rect 9585 11033 9597 11067
rect 9631 11064 9643 11067
rect 9950 11064 9956 11076
rect 9631 11036 9956 11064
rect 9631 11033 9643 11036
rect 9585 11027 9643 11033
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 10520 11064 10548 11092
rect 11624 11064 11652 11095
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 11793 11135 11851 11141
rect 11793 11132 11805 11135
rect 11756 11104 11805 11132
rect 11756 11092 11762 11104
rect 11793 11101 11805 11104
rect 11839 11101 11851 11135
rect 11900 11132 11928 11160
rect 11977 11135 12035 11141
rect 11977 11132 11989 11135
rect 11900 11104 11989 11132
rect 11793 11095 11851 11101
rect 11977 11101 11989 11104
rect 12023 11101 12035 11135
rect 11977 11095 12035 11101
rect 12250 11092 12256 11144
rect 12308 11092 12314 11144
rect 12360 11132 12388 11172
rect 13648 11172 14841 11200
rect 12509 11135 12567 11141
rect 12509 11132 12521 11135
rect 12360 11104 12521 11132
rect 12509 11101 12521 11104
rect 12555 11101 12567 11135
rect 12509 11095 12567 11101
rect 10520 11036 11652 11064
rect 11885 11067 11943 11073
rect 11885 11033 11897 11067
rect 11931 11064 11943 11067
rect 13648 11064 13676 11172
rect 14829 11169 14841 11172
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 14918 11160 14924 11212
rect 14976 11160 14982 11212
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11132 14795 11135
rect 15488 11132 15516 11296
rect 15746 11228 15752 11280
rect 15804 11228 15810 11280
rect 14783 11104 15516 11132
rect 14783 11101 14795 11104
rect 14737 11095 14795 11101
rect 11931 11036 13676 11064
rect 15381 11067 15439 11073
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 15381 11033 15393 11067
rect 15427 11064 15439 11067
rect 16114 11064 16120 11076
rect 15427 11036 16120 11064
rect 15427 11033 15439 11036
rect 15381 11027 15439 11033
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 6362 10996 6368 11008
rect 4632 10968 6368 10996
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 7006 10956 7012 11008
rect 7064 10956 7070 11008
rect 7466 10956 7472 11008
rect 7524 10956 7530 11008
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 8589 10999 8647 11005
rect 8589 10996 8601 10999
rect 8536 10968 8601 10996
rect 8536 10956 8542 10968
rect 8589 10965 8601 10968
rect 8635 10965 8647 10999
rect 8589 10959 8647 10965
rect 1104 10906 16811 10928
rect 1104 10854 4836 10906
rect 4888 10854 4900 10906
rect 4952 10854 4964 10906
rect 5016 10854 5028 10906
rect 5080 10854 5092 10906
rect 5144 10854 8723 10906
rect 8775 10854 8787 10906
rect 8839 10854 8851 10906
rect 8903 10854 8915 10906
rect 8967 10854 8979 10906
rect 9031 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 16497 10906
rect 16549 10854 16561 10906
rect 16613 10854 16625 10906
rect 16677 10854 16689 10906
rect 16741 10854 16753 10906
rect 16805 10854 16811 10906
rect 1104 10832 16811 10854
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 2869 10795 2927 10801
rect 2869 10792 2881 10795
rect 2832 10764 2881 10792
rect 2832 10752 2838 10764
rect 2869 10761 2881 10764
rect 2915 10761 2927 10795
rect 2869 10755 2927 10761
rect 3237 10795 3295 10801
rect 3237 10761 3249 10795
rect 3283 10792 3295 10795
rect 3326 10792 3332 10804
rect 3283 10764 3332 10792
rect 3283 10761 3295 10764
rect 3237 10755 3295 10761
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 4154 10752 4160 10804
rect 4212 10752 4218 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 4985 10795 5043 10801
rect 4985 10792 4997 10795
rect 4764 10764 4997 10792
rect 4764 10752 4770 10764
rect 4985 10761 4997 10764
rect 5031 10761 5043 10795
rect 4985 10755 5043 10761
rect 5810 10752 5816 10804
rect 5868 10752 5874 10804
rect 6086 10752 6092 10804
rect 6144 10752 6150 10804
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 6696 10764 6837 10792
rect 6696 10752 6702 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 7006 10752 7012 10804
rect 7064 10752 7070 10804
rect 7466 10752 7472 10804
rect 7524 10752 7530 10804
rect 8478 10752 8484 10804
rect 8536 10752 8542 10804
rect 8941 10795 8999 10801
rect 8941 10761 8953 10795
rect 8987 10792 8999 10795
rect 9398 10792 9404 10804
rect 8987 10764 9404 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 9585 10795 9643 10801
rect 9585 10792 9597 10795
rect 9548 10764 9597 10792
rect 9548 10752 9554 10764
rect 9585 10761 9597 10764
rect 9631 10761 9643 10795
rect 9585 10755 9643 10761
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 9824 10764 10977 10792
rect 9824 10752 9830 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 12066 10792 12072 10804
rect 11756 10764 12072 10792
rect 11756 10752 11762 10764
rect 12066 10752 12072 10764
rect 12124 10752 12130 10804
rect 14274 10752 14280 10804
rect 14332 10752 14338 10804
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10792 14979 10795
rect 15010 10792 15016 10804
rect 14967 10764 15016 10792
rect 14967 10761 14979 10764
rect 14921 10755 14979 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 15194 10752 15200 10804
rect 15252 10752 15258 10804
rect 1670 10733 1676 10736
rect 1664 10724 1676 10733
rect 1631 10696 1676 10724
rect 1664 10687 1676 10696
rect 1670 10684 1676 10687
rect 1728 10684 1734 10736
rect 4172 10724 4200 10752
rect 6104 10724 6132 10752
rect 3344 10696 4200 10724
rect 5184 10696 6132 10724
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10656 1455 10659
rect 2038 10656 2044 10668
rect 1443 10628 2044 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 3344 10665 3372 10696
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 3694 10616 3700 10668
rect 3752 10616 3758 10668
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 5184 10665 5212 10696
rect 7024 10665 7052 10752
rect 8294 10684 8300 10736
rect 8352 10684 8358 10736
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3936 10628 4077 10656
rect 3936 10616 3942 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10656 8263 10659
rect 8312 10656 8340 10684
rect 8251 10628 8340 10656
rect 8496 10656 8524 10752
rect 9674 10724 9680 10736
rect 9232 10696 9680 10724
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 8496 10628 8769 10656
rect 8251 10625 8263 10628
rect 8205 10619 8263 10625
rect 8757 10625 8769 10628
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 3513 10591 3571 10597
rect 3513 10557 3525 10591
rect 3559 10588 3571 10591
rect 3559 10560 3648 10588
rect 3559 10557 3571 10560
rect 3513 10551 3571 10557
rect 2777 10455 2835 10461
rect 2777 10421 2789 10455
rect 2823 10452 2835 10455
rect 3510 10452 3516 10464
rect 2823 10424 3516 10452
rect 2823 10421 2835 10424
rect 2777 10415 2835 10421
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 3620 10452 3648 10560
rect 3712 10520 3740 10616
rect 4338 10548 4344 10600
rect 4396 10548 4402 10600
rect 5350 10548 5356 10600
rect 5408 10588 5414 10600
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 5408 10560 5457 10588
rect 5408 10548 5414 10560
rect 5445 10557 5457 10560
rect 5491 10557 5503 10591
rect 5445 10551 5503 10557
rect 5644 10520 5672 10619
rect 7101 10591 7159 10597
rect 7101 10557 7113 10591
rect 7147 10588 7159 10591
rect 7190 10588 7196 10600
rect 7147 10560 7196 10588
rect 7147 10557 7159 10560
rect 7101 10551 7159 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7300 10520 7328 10619
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 8110 10588 8116 10600
rect 8067 10560 8116 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8570 10588 8576 10600
rect 8435 10560 8576 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 8864 10588 8892 10619
rect 9122 10588 9128 10600
rect 8864 10560 9128 10588
rect 8294 10520 8300 10532
rect 3712 10492 8300 10520
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 8864 10520 8892 10560
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9232 10597 9260 10696
rect 9600 10665 9628 10696
rect 9674 10684 9680 10696
rect 9732 10724 9738 10736
rect 10505 10727 10563 10733
rect 10505 10724 10517 10727
rect 9732 10696 10517 10724
rect 9732 10684 9738 10696
rect 10505 10693 10517 10696
rect 10551 10724 10563 10727
rect 10594 10724 10600 10736
rect 10551 10696 10600 10724
rect 10551 10693 10563 10696
rect 10505 10687 10563 10693
rect 10594 10684 10600 10696
rect 10652 10684 10658 10736
rect 14292 10724 14320 10752
rect 14292 10696 14872 10724
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 10134 10656 10140 10668
rect 9585 10619 9643 10625
rect 9692 10628 10140 10656
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 9416 10588 9444 10619
rect 9490 10588 9496 10600
rect 9416 10560 9496 10588
rect 9217 10551 9275 10557
rect 9490 10548 9496 10560
rect 9548 10588 9554 10600
rect 9692 10588 9720 10628
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 11054 10656 11060 10668
rect 10428 10628 11060 10656
rect 9548 10560 9720 10588
rect 9548 10548 9554 10560
rect 9766 10548 9772 10600
rect 9824 10548 9830 10600
rect 10428 10520 10456 10628
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11241 10659 11299 10665
rect 11241 10625 11253 10659
rect 11287 10656 11299 10659
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11287 10628 11529 10656
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 13906 10616 13912 10668
rect 13964 10656 13970 10668
rect 14274 10656 14280 10668
rect 13964 10628 14280 10656
rect 13964 10616 13970 10628
rect 14274 10616 14280 10628
rect 14332 10656 14338 10668
rect 14844 10665 14872 10696
rect 14461 10659 14519 10665
rect 14461 10656 14473 10659
rect 14332 10628 14473 10656
rect 14332 10616 14338 10628
rect 14461 10625 14473 10628
rect 14507 10625 14519 10659
rect 14461 10619 14519 10625
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 15010 10656 15016 10668
rect 14875 10628 15016 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 15212 10656 15240 10752
rect 15289 10659 15347 10665
rect 15289 10656 15301 10659
rect 15212 10628 15301 10656
rect 15289 10625 15301 10628
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 8404 10492 8892 10520
rect 9048 10492 10456 10520
rect 10505 10523 10563 10529
rect 8404 10464 8432 10492
rect 4062 10452 4068 10464
rect 3620 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 8386 10412 8392 10464
rect 8444 10412 8450 10464
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10452 8539 10455
rect 9048 10452 9076 10492
rect 10505 10489 10517 10523
rect 10551 10489 10563 10523
rect 10505 10483 10563 10489
rect 8527 10424 9076 10452
rect 9125 10455 9183 10461
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 9125 10421 9137 10455
rect 9171 10452 9183 10455
rect 9766 10452 9772 10464
rect 9171 10424 9772 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 10520 10452 10548 10483
rect 10192 10424 10548 10452
rect 10192 10412 10198 10424
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 13780 10424 14657 10452
rect 13780 10412 13786 10424
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 14645 10415 14703 10421
rect 15102 10412 15108 10464
rect 15160 10412 15166 10464
rect 1104 10362 16652 10384
rect 1104 10310 2893 10362
rect 2945 10310 2957 10362
rect 3009 10310 3021 10362
rect 3073 10310 3085 10362
rect 3137 10310 3149 10362
rect 3201 10310 6780 10362
rect 6832 10310 6844 10362
rect 6896 10310 6908 10362
rect 6960 10310 6972 10362
rect 7024 10310 7036 10362
rect 7088 10310 10667 10362
rect 10719 10310 10731 10362
rect 10783 10310 10795 10362
rect 10847 10310 10859 10362
rect 10911 10310 10923 10362
rect 10975 10310 14554 10362
rect 14606 10310 14618 10362
rect 14670 10310 14682 10362
rect 14734 10310 14746 10362
rect 14798 10310 14810 10362
rect 14862 10310 16652 10362
rect 1104 10288 16652 10310
rect 5534 10208 5540 10260
rect 5592 10208 5598 10260
rect 5644 10220 7328 10248
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 5644 10180 5672 10220
rect 5408 10152 5672 10180
rect 7300 10180 7328 10220
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 9398 10248 9404 10260
rect 8352 10220 9404 10248
rect 8352 10208 8358 10220
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 9674 10208 9680 10260
rect 9732 10208 9738 10260
rect 9950 10208 9956 10260
rect 10008 10208 10014 10260
rect 11146 10208 11152 10260
rect 11204 10248 11210 10260
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 11204 10220 11437 10248
rect 11204 10208 11210 10220
rect 11425 10217 11437 10220
rect 11471 10248 11483 10251
rect 11882 10248 11888 10260
rect 11471 10220 11888 10248
rect 11471 10217 11483 10220
rect 11425 10211 11483 10217
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 13906 10248 13912 10260
rect 12176 10220 13912 10248
rect 9122 10180 9128 10192
rect 7300 10152 9128 10180
rect 5408 10140 5414 10152
rect 9122 10140 9128 10152
rect 9180 10180 9186 10192
rect 9180 10152 11376 10180
rect 9180 10140 9186 10152
rect 2038 10072 2044 10124
rect 2096 10112 2102 10124
rect 3789 10115 3847 10121
rect 3789 10112 3801 10115
rect 2096 10084 3801 10112
rect 2096 10072 2102 10084
rect 3789 10081 3801 10084
rect 3835 10112 3847 10115
rect 6362 10112 6368 10124
rect 3835 10084 6368 10112
rect 3835 10081 3847 10084
rect 3789 10075 3847 10081
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 9950 10112 9956 10124
rect 9723 10084 9956 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 9950 10072 9956 10084
rect 10008 10112 10014 10124
rect 10318 10112 10324 10124
rect 10008 10084 10324 10112
rect 10008 10072 10014 10084
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 3602 10004 3608 10056
rect 3660 10004 3666 10056
rect 5626 10004 5632 10056
rect 5684 10044 5690 10056
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5684 10016 5733 10044
rect 5684 10004 5690 10016
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 9585 10047 9643 10053
rect 9585 10013 9597 10047
rect 9631 10013 9643 10047
rect 9585 10007 9643 10013
rect 4065 9979 4123 9985
rect 4065 9976 4077 9979
rect 3436 9948 4077 9976
rect 3436 9917 3464 9948
rect 4065 9945 4077 9948
rect 4111 9945 4123 9979
rect 4065 9939 4123 9945
rect 4522 9936 4528 9988
rect 4580 9936 4586 9988
rect 5736 9976 5764 10007
rect 6632 9979 6690 9985
rect 5736 9948 6592 9976
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9877 3479 9911
rect 3421 9871 3479 9877
rect 5997 9911 6055 9917
rect 5997 9877 6009 9911
rect 6043 9908 6055 9911
rect 6178 9908 6184 9920
rect 6043 9880 6184 9908
rect 6043 9877 6055 9880
rect 5997 9871 6055 9877
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 6564 9908 6592 9948
rect 6632 9945 6644 9979
rect 6678 9976 6690 9979
rect 6914 9976 6920 9988
rect 6678 9948 6920 9976
rect 6678 9945 6690 9948
rect 6632 9939 6690 9945
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 9125 9979 9183 9985
rect 9125 9945 9137 9979
rect 9171 9976 9183 9979
rect 9306 9976 9312 9988
rect 9171 9948 9312 9976
rect 9171 9945 9183 9948
rect 9125 9939 9183 9945
rect 7745 9911 7803 9917
rect 7745 9908 7757 9911
rect 6564 9880 7757 9908
rect 7745 9877 7757 9880
rect 7791 9908 7803 9911
rect 9140 9908 9168 9939
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 9600 9976 9628 10007
rect 11238 10004 11244 10056
rect 11296 10004 11302 10056
rect 11348 10044 11376 10152
rect 11900 10112 11928 10208
rect 11900 10084 12020 10112
rect 11885 10047 11943 10053
rect 11885 10044 11897 10047
rect 11348 10016 11897 10044
rect 11885 10013 11897 10016
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 9766 9976 9772 9988
rect 9600 9948 9772 9976
rect 9600 9920 9628 9948
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 7791 9880 9168 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 9398 9868 9404 9920
rect 9456 9868 9462 9920
rect 9582 9868 9588 9920
rect 9640 9868 9646 9920
rect 11992 9908 12020 10084
rect 12066 10004 12072 10056
rect 12124 10004 12130 10056
rect 12176 10053 12204 10220
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 12492 10084 12541 10112
rect 12492 10072 12498 10084
rect 12529 10081 12541 10084
rect 12575 10081 12587 10115
rect 12529 10075 12587 10081
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10112 14795 10115
rect 15102 10112 15108 10124
rect 14783 10084 15108 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12544 10044 12572 10075
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 13722 10044 13728 10056
rect 12544 10016 13728 10044
rect 12253 10007 12311 10013
rect 12268 9976 12296 10007
rect 13722 10004 13728 10016
rect 13780 10044 13786 10056
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 13780 10016 14473 10044
rect 13780 10004 13786 10016
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 12774 9979 12832 9985
rect 12774 9976 12786 9979
rect 12176 9948 12296 9976
rect 12452 9948 12786 9976
rect 12176 9908 12204 9948
rect 12452 9917 12480 9948
rect 12774 9945 12786 9948
rect 12820 9945 12832 9979
rect 12774 9939 12832 9945
rect 15378 9936 15384 9988
rect 15436 9936 15442 9988
rect 11992 9880 12204 9908
rect 12437 9911 12495 9917
rect 12437 9877 12449 9911
rect 12483 9877 12495 9911
rect 12437 9871 12495 9877
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 16209 9911 16267 9917
rect 16209 9908 16221 9911
rect 14608 9880 16221 9908
rect 14608 9868 14614 9880
rect 16209 9877 16221 9880
rect 16255 9877 16267 9911
rect 16209 9871 16267 9877
rect 1104 9818 16811 9840
rect 1104 9766 4836 9818
rect 4888 9766 4900 9818
rect 4952 9766 4964 9818
rect 5016 9766 5028 9818
rect 5080 9766 5092 9818
rect 5144 9766 8723 9818
rect 8775 9766 8787 9818
rect 8839 9766 8851 9818
rect 8903 9766 8915 9818
rect 8967 9766 8979 9818
rect 9031 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 16497 9818
rect 16549 9766 16561 9818
rect 16613 9766 16625 9818
rect 16677 9766 16689 9818
rect 16741 9766 16753 9818
rect 16805 9766 16811 9818
rect 1104 9744 16811 9766
rect 3513 9707 3571 9713
rect 3513 9673 3525 9707
rect 3559 9704 3571 9707
rect 3602 9704 3608 9716
rect 3559 9676 3608 9704
rect 3559 9673 3571 9676
rect 3513 9667 3571 9673
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 4522 9664 4528 9716
rect 4580 9664 4586 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6641 9707 6699 9713
rect 6641 9704 6653 9707
rect 6420 9676 6653 9704
rect 6420 9664 6426 9676
rect 6641 9673 6653 9676
rect 6687 9673 6699 9707
rect 6641 9667 6699 9673
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 9674 9664 9680 9716
rect 9732 9664 9738 9716
rect 12066 9704 12072 9716
rect 10980 9676 12072 9704
rect 4338 9596 4344 9648
rect 4396 9636 4402 9648
rect 4396 9608 4476 9636
rect 4396 9596 4402 9608
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9568 1455 9571
rect 1486 9568 1492 9580
rect 1443 9540 1492 9568
rect 1443 9537 1455 9540
rect 1397 9531 1455 9537
rect 1486 9528 1492 9540
rect 1544 9528 1550 9580
rect 1670 9577 1676 9580
rect 1664 9531 1676 9577
rect 1670 9528 1676 9531
rect 1728 9528 1734 9580
rect 3878 9528 3884 9580
rect 3936 9528 3942 9580
rect 4448 9577 4476 9608
rect 6178 9596 6184 9648
rect 6236 9636 6242 9648
rect 7837 9639 7895 9645
rect 7837 9636 7849 9639
rect 6236 9608 7849 9636
rect 6236 9596 6242 9608
rect 7837 9605 7849 9608
rect 7883 9605 7895 9639
rect 7837 9599 7895 9605
rect 7929 9639 7987 9645
rect 7929 9605 7941 9639
rect 7975 9636 7987 9639
rect 8389 9639 8447 9645
rect 8389 9636 8401 9639
rect 7975 9608 8401 9636
rect 7975 9605 7987 9608
rect 7929 9599 7987 9605
rect 8389 9605 8401 9608
rect 8435 9605 8447 9639
rect 8389 9599 8447 9605
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9500 4123 9503
rect 4154 9500 4160 9512
rect 4111 9472 4160 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 2774 9392 2780 9444
rect 2832 9432 2838 9444
rect 3988 9432 4016 9463
rect 4154 9460 4160 9472
rect 4212 9500 4218 9512
rect 6196 9500 6224 9596
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9568 6515 9571
rect 6546 9568 6552 9580
rect 6503 9540 6552 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9568 7159 9571
rect 7147 9540 7512 9568
rect 7147 9537 7159 9540
rect 7101 9531 7159 9537
rect 4212 9472 6224 9500
rect 4212 9460 4218 9472
rect 7484 9441 7512 9540
rect 8294 9528 8300 9580
rect 8352 9528 8358 9580
rect 8478 9528 8484 9580
rect 8536 9528 8542 9580
rect 8846 9528 8852 9580
rect 8904 9568 8910 9580
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 8904 9540 8953 9568
rect 8904 9528 8910 9540
rect 8941 9537 8953 9540
rect 8987 9568 8999 9571
rect 9692 9568 9720 9664
rect 10980 9645 11008 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 13906 9664 13912 9716
rect 13964 9664 13970 9716
rect 14550 9664 14556 9716
rect 14608 9664 14614 9716
rect 15378 9664 15384 9716
rect 15436 9664 15442 9716
rect 10965 9639 11023 9645
rect 10965 9605 10977 9639
rect 11011 9605 11023 9639
rect 13924 9636 13952 9664
rect 14645 9639 14703 9645
rect 14645 9636 14657 9639
rect 10965 9599 11023 9605
rect 11072 9608 12434 9636
rect 13924 9608 14657 9636
rect 8987 9540 9720 9568
rect 10137 9571 10195 9577
rect 8987 9537 8999 9540
rect 8941 9531 8999 9537
rect 10137 9537 10149 9571
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9500 8171 9503
rect 8570 9500 8576 9512
rect 8159 9472 8576 9500
rect 8159 9469 8171 9472
rect 8113 9463 8171 9469
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9490 9500 9496 9512
rect 9263 9472 9496 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 10152 9500 10180 9531
rect 10410 9528 10416 9580
rect 10468 9568 10474 9580
rect 11072 9577 11100 9608
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10468 9540 10793 9568
rect 10468 9528 10474 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 11146 9528 11152 9580
rect 11204 9528 11210 9580
rect 11773 9571 11831 9577
rect 11773 9568 11785 9571
rect 11348 9540 11785 9568
rect 10318 9500 10324 9512
rect 10152 9472 10324 9500
rect 2832 9404 4016 9432
rect 7469 9435 7527 9441
rect 2832 9392 2838 9404
rect 7469 9401 7481 9435
rect 7515 9401 7527 9435
rect 9582 9432 9588 9444
rect 7469 9395 7527 9401
rect 9324 9404 9588 9432
rect 9324 9376 9352 9404
rect 9582 9392 9588 9404
rect 9640 9432 9646 9444
rect 10152 9432 10180 9472
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 11348 9441 11376 9540
rect 11773 9537 11785 9540
rect 11819 9537 11831 9571
rect 12406 9568 12434 9608
rect 14645 9605 14657 9608
rect 14691 9605 14703 9639
rect 14645 9599 14703 9605
rect 15010 9596 15016 9648
rect 15068 9636 15074 9648
rect 15068 9608 15332 9636
rect 15068 9596 15074 9608
rect 15304 9577 15332 9608
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 12406 9540 12848 9568
rect 11773 9531 11831 9537
rect 11517 9503 11575 9509
rect 11517 9469 11529 9503
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 9640 9404 10180 9432
rect 11333 9435 11391 9441
rect 9640 9392 9646 9404
rect 11333 9401 11345 9435
rect 11379 9401 11391 9435
rect 11333 9395 11391 9401
rect 9306 9324 9312 9376
rect 9364 9324 9370 9376
rect 9490 9324 9496 9376
rect 9548 9324 9554 9376
rect 10226 9324 10232 9376
rect 10284 9324 10290 9376
rect 11532 9364 11560 9463
rect 12820 9432 12848 9540
rect 14200 9540 15209 9568
rect 12894 9432 12900 9444
rect 12820 9404 12900 9432
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 14200 9441 14228 9540
rect 15197 9537 15209 9540
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 15289 9571 15347 9577
rect 15289 9537 15301 9571
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 16298 9528 16304 9580
rect 16356 9528 16362 9580
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 14918 9500 14924 9512
rect 14875 9472 14924 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 14185 9435 14243 9441
rect 14185 9401 14197 9435
rect 14231 9401 14243 9435
rect 14185 9395 14243 9401
rect 11882 9364 11888 9376
rect 11532 9336 11888 9364
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 15010 9324 15016 9376
rect 15068 9324 15074 9376
rect 1104 9274 16652 9296
rect 1104 9222 2893 9274
rect 2945 9222 2957 9274
rect 3009 9222 3021 9274
rect 3073 9222 3085 9274
rect 3137 9222 3149 9274
rect 3201 9222 6780 9274
rect 6832 9222 6844 9274
rect 6896 9222 6908 9274
rect 6960 9222 6972 9274
rect 7024 9222 7036 9274
rect 7088 9222 10667 9274
rect 10719 9222 10731 9274
rect 10783 9222 10795 9274
rect 10847 9222 10859 9274
rect 10911 9222 10923 9274
rect 10975 9222 14554 9274
rect 14606 9222 14618 9274
rect 14670 9222 14682 9274
rect 14734 9222 14746 9274
rect 14798 9222 14810 9274
rect 14862 9222 16652 9274
rect 1104 9200 16652 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 1670 9160 1676 9172
rect 1627 9132 1676 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 2774 9160 2780 9172
rect 2746 9120 2780 9160
rect 2832 9120 2838 9172
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8478 9160 8484 9172
rect 7975 9132 8484 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 8757 9163 8815 9169
rect 8757 9129 8769 9163
rect 8803 9160 8815 9163
rect 9306 9160 9312 9172
rect 8803 9132 9312 9160
rect 8803 9129 8815 9132
rect 8757 9123 8815 9129
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 9490 9120 9496 9172
rect 9548 9120 9554 9172
rect 9858 9120 9864 9172
rect 9916 9160 9922 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 9916 9132 10241 9160
rect 9916 9120 9922 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 11149 9163 11207 9169
rect 11149 9129 11161 9163
rect 11195 9129 11207 9163
rect 11149 9123 11207 9129
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 9024 2559 9027
rect 2590 9024 2596 9036
rect 2547 8996 2596 9024
rect 2547 8993 2559 8996
rect 2501 8987 2559 8993
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 2225 8959 2283 8965
rect 1811 8928 1900 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 1872 8829 1900 8928
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2746 8956 2774 9120
rect 8294 9052 8300 9104
rect 8352 9052 8358 9104
rect 4338 9024 4344 9036
rect 3896 8996 4344 9024
rect 3896 8965 3924 8996
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 5442 8984 5448 9036
rect 5500 8984 5506 9036
rect 8018 9024 8024 9036
rect 7852 8996 8024 9024
rect 2271 8928 2774 8956
rect 3881 8959 3939 8965
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 3881 8925 3893 8959
rect 3927 8925 3939 8959
rect 3881 8919 3939 8925
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 7852 8965 7880 8996
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8925 7895 8959
rect 7837 8919 7895 8925
rect 5644 8888 5672 8919
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 8312 8888 8340 9052
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 8536 8996 8953 9024
rect 8536 8984 8542 8996
rect 8941 8993 8953 8996
rect 8987 9024 8999 9027
rect 9508 9024 9536 9120
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 10689 9095 10747 9101
rect 10689 9092 10701 9095
rect 9732 9064 10701 9092
rect 9732 9052 9738 9064
rect 10689 9061 10701 9064
rect 10735 9061 10747 9095
rect 10689 9055 10747 9061
rect 10873 9095 10931 9101
rect 10873 9061 10885 9095
rect 10919 9092 10931 9095
rect 11164 9092 11192 9123
rect 11238 9120 11244 9172
rect 11296 9160 11302 9172
rect 11425 9163 11483 9169
rect 11425 9160 11437 9163
rect 11296 9132 11437 9160
rect 11296 9120 11302 9132
rect 11425 9129 11437 9132
rect 11471 9129 11483 9163
rect 11425 9123 11483 9129
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9129 11759 9163
rect 11701 9123 11759 9129
rect 11716 9092 11744 9123
rect 12894 9120 12900 9172
rect 12952 9120 12958 9172
rect 14918 9160 14924 9172
rect 14108 9132 14924 9160
rect 10919 9064 11744 9092
rect 10919 9061 10931 9064
rect 10873 9055 10931 9061
rect 10134 9024 10140 9036
rect 8987 8996 9536 9024
rect 9784 8996 10140 9024
rect 8987 8993 8999 8996
rect 8941 8987 8999 8993
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 8846 8956 8852 8968
rect 8619 8928 8852 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9140 8888 9168 8919
rect 9214 8916 9220 8968
rect 9272 8956 9278 8968
rect 9784 8965 9812 8996
rect 10134 8984 10140 8996
rect 10192 9024 10198 9036
rect 10413 9027 10471 9033
rect 10413 9024 10425 9027
rect 10192 8996 10425 9024
rect 10192 8984 10198 8996
rect 10413 8993 10425 8996
rect 10459 8993 10471 9027
rect 10413 8987 10471 8993
rect 11054 8984 11060 9036
rect 11112 8984 11118 9036
rect 12912 9024 12940 9120
rect 13081 9027 13139 9033
rect 13081 9024 13093 9027
rect 12912 8996 13093 9024
rect 13081 8993 13093 8996
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 14108 9024 14136 9132
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 13311 8996 14136 9024
rect 14369 9027 14427 9033
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 14369 8993 14381 9027
rect 14415 9024 14427 9027
rect 15010 9024 15016 9036
rect 14415 8996 15016 9024
rect 14415 8993 14427 8996
rect 14369 8987 14427 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 15102 8984 15108 9036
rect 15160 9024 15166 9036
rect 15160 8996 15976 9024
rect 15160 8984 15166 8996
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 9272 8928 9321 8956
rect 9272 8916 9278 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 10226 8956 10232 8968
rect 9907 8928 10232 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 10226 8916 10232 8928
rect 10284 8956 10290 8968
rect 10965 8959 11023 8965
rect 10284 8928 10548 8956
rect 10284 8916 10290 8928
rect 5644 8860 8156 8888
rect 8128 8832 8156 8860
rect 8312 8860 9168 8888
rect 10520 8888 10548 8928
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 11072 8956 11100 8984
rect 11011 8928 11652 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11514 8888 11520 8900
rect 10520 8860 11520 8888
rect 1857 8823 1915 8829
rect 1857 8789 1869 8823
rect 1903 8789 1915 8823
rect 1857 8783 1915 8789
rect 2314 8780 2320 8832
rect 2372 8780 2378 8832
rect 3970 8780 3976 8832
rect 4028 8780 4034 8832
rect 5166 8780 5172 8832
rect 5224 8780 5230 8832
rect 5810 8780 5816 8832
rect 5868 8780 5874 8832
rect 8110 8780 8116 8832
rect 8168 8780 8174 8832
rect 8312 8820 8340 8860
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 11624 8888 11652 8928
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 15948 8965 15976 8996
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13964 8928 14105 8956
rect 13964 8916 13970 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8925 15991 8959
rect 15933 8919 15991 8925
rect 11717 8891 11775 8897
rect 11717 8888 11729 8891
rect 11624 8860 11729 8888
rect 11717 8857 11729 8860
rect 11763 8857 11775 8891
rect 11717 8851 11775 8857
rect 12989 8891 13047 8897
rect 12989 8857 13001 8891
rect 13035 8888 13047 8891
rect 16025 8891 16083 8897
rect 16025 8888 16037 8891
rect 13035 8860 14320 8888
rect 15594 8860 16037 8888
rect 13035 8857 13047 8860
rect 12989 8851 13047 8857
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8312 8792 8401 8820
rect 8389 8789 8401 8792
rect 8435 8820 8447 8823
rect 8570 8820 8576 8832
rect 8435 8792 8576 8820
rect 8435 8789 8447 8792
rect 8389 8783 8447 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 11882 8780 11888 8832
rect 11940 8780 11946 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 12621 8823 12679 8829
rect 12621 8820 12633 8823
rect 12584 8792 12633 8820
rect 12584 8780 12590 8792
rect 12621 8789 12633 8792
rect 12667 8789 12679 8823
rect 14292 8820 14320 8860
rect 16025 8857 16037 8860
rect 16071 8857 16083 8891
rect 16025 8851 16083 8857
rect 15841 8823 15899 8829
rect 15841 8820 15853 8823
rect 14292 8792 15853 8820
rect 12621 8783 12679 8789
rect 15841 8789 15853 8792
rect 15887 8789 15899 8823
rect 15841 8783 15899 8789
rect 1104 8730 16811 8752
rect 1104 8678 4836 8730
rect 4888 8678 4900 8730
rect 4952 8678 4964 8730
rect 5016 8678 5028 8730
rect 5080 8678 5092 8730
rect 5144 8678 8723 8730
rect 8775 8678 8787 8730
rect 8839 8678 8851 8730
rect 8903 8678 8915 8730
rect 8967 8678 8979 8730
rect 9031 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 16497 8730
rect 16549 8678 16561 8730
rect 16613 8678 16625 8730
rect 16677 8678 16689 8730
rect 16741 8678 16753 8730
rect 16805 8678 16811 8730
rect 1104 8656 16811 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2409 8619 2467 8625
rect 2409 8616 2421 8619
rect 2372 8588 2421 8616
rect 2372 8576 2378 8588
rect 2409 8585 2421 8588
rect 2455 8585 2467 8619
rect 2409 8579 2467 8585
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 3936 8588 4353 8616
rect 3936 8576 3942 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 4341 8579 4399 8585
rect 5166 8576 5172 8628
rect 5224 8576 5230 8628
rect 8478 8576 8484 8628
rect 8536 8576 8542 8628
rect 8570 8576 8576 8628
rect 8628 8576 8634 8628
rect 11514 8576 11520 8628
rect 11572 8576 11578 8628
rect 12526 8576 12532 8628
rect 12584 8576 12590 8628
rect 1486 8508 1492 8560
rect 1544 8548 1550 8560
rect 1544 8520 2636 8548
rect 1544 8508 1550 8520
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8480 2283 8483
rect 2498 8480 2504 8492
rect 2271 8452 2504 8480
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 2608 8489 2636 8520
rect 2774 8508 2780 8560
rect 2832 8548 2838 8560
rect 2869 8551 2927 8557
rect 2869 8548 2881 8551
rect 2832 8520 2881 8548
rect 2832 8508 2838 8520
rect 2869 8517 2881 8520
rect 2915 8517 2927 8551
rect 2869 8511 2927 8517
rect 5068 8551 5126 8557
rect 5068 8517 5080 8551
rect 5114 8548 5126 8551
rect 5184 8548 5212 8576
rect 7190 8548 7196 8560
rect 5114 8520 5212 8548
rect 6932 8520 7196 8548
rect 5114 8517 5126 8520
rect 5068 8511 5126 8517
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 3970 8440 3976 8492
rect 4028 8440 4034 8492
rect 6932 8480 6960 8520
rect 7190 8508 7196 8520
rect 7248 8508 7254 8560
rect 4448 8452 6960 8480
rect 7009 8483 7067 8489
rect 2041 8415 2099 8421
rect 2041 8381 2053 8415
rect 2087 8381 2099 8415
rect 4448 8412 4476 8452
rect 7009 8449 7021 8483
rect 7055 8480 7067 8483
rect 7098 8480 7104 8492
rect 7055 8452 7104 8480
rect 7055 8449 7067 8452
rect 7009 8443 7067 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 2041 8375 2099 8381
rect 2700 8384 4476 8412
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2056 8344 2084 8375
rect 2700 8344 2728 8384
rect 4522 8372 4528 8424
rect 4580 8412 4586 8424
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 4580 8384 4813 8412
rect 4580 8372 4586 8384
rect 4801 8381 4813 8384
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 1627 8316 2728 8344
rect 7208 8344 7236 8508
rect 8496 8489 8524 8576
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 8588 8480 8616 8576
rect 11532 8548 11560 8576
rect 10704 8520 11560 8548
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 8588 8452 8677 8480
rect 8481 8443 8539 8449
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 9214 8480 9220 8492
rect 8895 8452 9220 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 9030 8412 9036 8424
rect 8260 8384 9036 8412
rect 8260 8372 8266 8384
rect 9030 8372 9036 8384
rect 9088 8412 9094 8424
rect 9324 8412 9352 8443
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 9674 8480 9680 8492
rect 9456 8452 9680 8480
rect 9456 8440 9462 8452
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 10704 8489 10732 8520
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 11054 8440 11060 8492
rect 11112 8440 11118 8492
rect 12544 8480 12572 8576
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12544 8452 12909 8480
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 10152 8412 10180 8440
rect 9088 8384 10180 8412
rect 9088 8372 9094 8384
rect 10318 8372 10324 8424
rect 10376 8412 10382 8424
rect 12434 8412 12440 8424
rect 10376 8384 12440 8412
rect 10376 8372 10382 8384
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 9674 8344 9680 8356
rect 7208 8316 9680 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 9674 8304 9680 8316
rect 9732 8344 9738 8356
rect 10410 8344 10416 8356
rect 9732 8316 10416 8344
rect 9732 8304 9738 8316
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 11790 8344 11796 8356
rect 11112 8316 11796 8344
rect 11112 8304 11118 8316
rect 11790 8304 11796 8316
rect 11848 8304 11854 8356
rect 6178 8236 6184 8288
rect 6236 8236 6242 8288
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6696 8248 6837 8276
rect 6696 8236 6702 8248
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 9769 8279 9827 8285
rect 9769 8276 9781 8279
rect 8536 8248 9781 8276
rect 8536 8236 8542 8248
rect 9769 8245 9781 8248
rect 9815 8245 9827 8279
rect 9769 8239 9827 8245
rect 12526 8236 12532 8288
rect 12584 8276 12590 8288
rect 12713 8279 12771 8285
rect 12713 8276 12725 8279
rect 12584 8248 12725 8276
rect 12584 8236 12590 8248
rect 12713 8245 12725 8248
rect 12759 8245 12771 8279
rect 12713 8239 12771 8245
rect 1104 8186 16652 8208
rect 1104 8134 2893 8186
rect 2945 8134 2957 8186
rect 3009 8134 3021 8186
rect 3073 8134 3085 8186
rect 3137 8134 3149 8186
rect 3201 8134 6780 8186
rect 6832 8134 6844 8186
rect 6896 8134 6908 8186
rect 6960 8134 6972 8186
rect 7024 8134 7036 8186
rect 7088 8134 10667 8186
rect 10719 8134 10731 8186
rect 10783 8134 10795 8186
rect 10847 8134 10859 8186
rect 10911 8134 10923 8186
rect 10975 8134 14554 8186
rect 14606 8134 14618 8186
rect 14670 8134 14682 8186
rect 14734 8134 14746 8186
rect 14798 8134 14810 8186
rect 14862 8134 16652 8186
rect 1104 8112 16652 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2832 8044 2973 8072
rect 2832 8032 2838 8044
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 5350 8032 5356 8084
rect 5408 8032 5414 8084
rect 9309 8075 9367 8081
rect 6472 8044 8524 8072
rect 2608 7976 6040 8004
rect 2608 7948 2636 7976
rect 2590 7896 2596 7948
rect 2648 7896 2654 7948
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4212 7908 4445 7936
rect 4212 7896 4218 7908
rect 4433 7905 4445 7908
rect 4479 7936 4491 7939
rect 5350 7936 5356 7948
rect 4479 7908 5356 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5810 7896 5816 7948
rect 5868 7896 5874 7948
rect 6012 7945 6040 7976
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7936 6055 7939
rect 6472 7936 6500 8044
rect 8496 8016 8524 8044
rect 9309 8041 9321 8075
rect 9355 8072 9367 8075
rect 9398 8072 9404 8084
rect 9355 8044 9404 8072
rect 9355 8041 9367 8044
rect 9309 8035 9367 8041
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10962 8072 10968 8084
rect 10008 8044 10968 8072
rect 10008 8032 10014 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11882 8032 11888 8084
rect 11940 8032 11946 8084
rect 8478 7964 8484 8016
rect 8536 7964 8542 8016
rect 6043 7908 6500 7936
rect 7929 7939 7987 7945
rect 6043 7905 6055 7908
rect 5997 7899 6055 7905
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 9968 7936 9996 8032
rect 11054 8004 11060 8016
rect 7975 7908 9996 7936
rect 10060 7976 11060 8004
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7868 3203 7871
rect 3191 7840 3832 7868
rect 3191 7837 3203 7840
rect 3145 7831 3203 7837
rect 3804 7741 3832 7840
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 6178 7868 6184 7880
rect 5776 7840 6184 7868
rect 5776 7828 5782 7840
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 6713 7871 6771 7877
rect 6713 7868 6725 7871
rect 6656 7840 6725 7868
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 4249 7803 4307 7809
rect 4249 7800 4261 7803
rect 4120 7772 4261 7800
rect 4120 7760 4126 7772
rect 4249 7769 4261 7772
rect 4295 7769 4307 7803
rect 4249 7763 4307 7769
rect 6656 7744 6684 7840
rect 6713 7837 6725 7840
rect 6759 7837 6771 7871
rect 6713 7831 6771 7837
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8941 7871 8999 7877
rect 8168 7840 8616 7868
rect 8168 7828 8174 7840
rect 8588 7800 8616 7840
rect 8941 7837 8953 7871
rect 8987 7868 8999 7871
rect 9030 7868 9036 7880
rect 8987 7840 9036 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9232 7840 9597 7868
rect 9232 7800 9260 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9674 7828 9680 7880
rect 9732 7828 9738 7880
rect 10060 7877 10088 7976
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 11900 7936 11928 8032
rect 10888 7908 11928 7936
rect 12437 7939 12495 7945
rect 10888 7877 10916 7908
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 12526 7936 12532 7948
rect 12483 7908 12532 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 14737 7939 14795 7945
rect 14737 7905 14749 7939
rect 14783 7936 14795 7939
rect 14918 7936 14924 7948
rect 14783 7908 14924 7936
rect 14783 7905 14795 7908
rect 14737 7899 14795 7905
rect 14918 7896 14924 7908
rect 14976 7896 14982 7948
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10873 7871 10931 7877
rect 10873 7837 10885 7871
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 11020 7840 11529 7868
rect 11020 7828 11026 7840
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 12032 7840 12173 7868
rect 12032 7828 12038 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14553 7871 14611 7877
rect 14553 7868 14565 7871
rect 13872 7840 14565 7868
rect 13872 7828 13878 7840
rect 14553 7837 14565 7840
rect 14599 7837 14611 7871
rect 14553 7831 14611 7837
rect 8588 7772 9260 7800
rect 8588 7744 8616 7772
rect 9306 7760 9312 7812
rect 9364 7809 9370 7812
rect 9364 7800 9376 7809
rect 9861 7803 9919 7809
rect 9364 7772 9409 7800
rect 9364 7763 9376 7772
rect 9861 7769 9873 7803
rect 9907 7769 9919 7803
rect 9861 7763 9919 7769
rect 9364 7760 9370 7763
rect 3789 7735 3847 7741
rect 3789 7701 3801 7735
rect 3835 7701 3847 7735
rect 3789 7695 3847 7701
rect 4154 7692 4160 7744
rect 4212 7692 4218 7744
rect 6638 7692 6644 7744
rect 6696 7692 6702 7744
rect 7374 7692 7380 7744
rect 7432 7732 7438 7744
rect 7837 7735 7895 7741
rect 7837 7732 7849 7735
rect 7432 7704 7849 7732
rect 7432 7692 7438 7704
rect 7837 7701 7849 7704
rect 7883 7701 7895 7735
rect 7837 7695 7895 7701
rect 8294 7692 8300 7744
rect 8352 7692 8358 7744
rect 8570 7692 8576 7744
rect 8628 7692 8634 7744
rect 9876 7732 9904 7763
rect 9950 7760 9956 7812
rect 10008 7760 10014 7812
rect 11701 7803 11759 7809
rect 11701 7800 11713 7803
rect 10060 7772 11713 7800
rect 10060 7732 10088 7772
rect 11164 7744 11192 7772
rect 11701 7769 11713 7772
rect 11747 7769 11759 7803
rect 11701 7763 11759 7769
rect 11793 7803 11851 7809
rect 11793 7769 11805 7803
rect 11839 7800 11851 7803
rect 13722 7800 13728 7812
rect 11839 7772 12434 7800
rect 13662 7772 13728 7800
rect 11839 7769 11851 7772
rect 11793 7763 11851 7769
rect 9876 7704 10088 7732
rect 10226 7692 10232 7744
rect 10284 7692 10290 7744
rect 11057 7735 11115 7741
rect 11057 7701 11069 7735
rect 11103 7732 11115 7735
rect 11146 7732 11152 7744
rect 11103 7704 11152 7732
rect 11103 7701 11115 7704
rect 11057 7695 11115 7701
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 12066 7692 12072 7744
rect 12124 7692 12130 7744
rect 12406 7732 12434 7772
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 13832 7732 13860 7828
rect 14461 7803 14519 7809
rect 14461 7800 14473 7803
rect 13924 7772 14473 7800
rect 13924 7741 13952 7772
rect 14461 7769 14473 7772
rect 14507 7769 14519 7803
rect 14461 7763 14519 7769
rect 12406 7704 13860 7732
rect 13909 7735 13967 7741
rect 13909 7701 13921 7735
rect 13955 7701 13967 7735
rect 13909 7695 13967 7701
rect 14090 7692 14096 7744
rect 14148 7692 14154 7744
rect 1104 7642 16811 7664
rect 1104 7590 4836 7642
rect 4888 7590 4900 7642
rect 4952 7590 4964 7642
rect 5016 7590 5028 7642
rect 5080 7590 5092 7642
rect 5144 7590 8723 7642
rect 8775 7590 8787 7642
rect 8839 7590 8851 7642
rect 8903 7590 8915 7642
rect 8967 7590 8979 7642
rect 9031 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 16497 7642
rect 16549 7590 16561 7642
rect 16613 7590 16625 7642
rect 16677 7590 16689 7642
rect 16741 7590 16753 7642
rect 16805 7590 16811 7642
rect 1104 7568 16811 7590
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 4062 7528 4068 7540
rect 2832 7500 4068 7528
rect 2832 7488 2838 7500
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 4212 7500 4905 7528
rect 4212 7488 4218 7500
rect 4893 7497 4905 7500
rect 4939 7497 4951 7531
rect 4893 7491 4951 7497
rect 5718 7488 5724 7540
rect 5776 7488 5782 7540
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 7098 7528 7104 7540
rect 7055 7500 7104 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 7374 7488 7380 7540
rect 7432 7488 7438 7540
rect 7469 7531 7527 7537
rect 7469 7497 7481 7531
rect 7515 7528 7527 7531
rect 8294 7528 8300 7540
rect 7515 7500 8300 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 10226 7488 10232 7540
rect 10284 7488 10290 7540
rect 12066 7488 12072 7540
rect 12124 7488 12130 7540
rect 13357 7531 13415 7537
rect 13357 7497 13369 7531
rect 13403 7497 13415 7531
rect 13357 7491 13415 7497
rect 5077 7463 5135 7469
rect 5077 7460 5089 7463
rect 1504 7432 2774 7460
rect 4646 7432 5089 7460
rect 1504 7404 1532 7432
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 1486 7392 1492 7404
rect 1443 7364 1492 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 1486 7352 1492 7364
rect 1544 7352 1550 7404
rect 1670 7401 1676 7404
rect 1664 7355 1676 7401
rect 1670 7352 1676 7355
rect 1728 7352 1734 7404
rect 2746 7324 2774 7432
rect 5077 7429 5089 7432
rect 5123 7429 5135 7463
rect 5077 7423 5135 7429
rect 8748 7463 8806 7469
rect 8748 7429 8760 7463
rect 8794 7460 8806 7463
rect 10244 7460 10272 7488
rect 8794 7432 10272 7460
rect 12084 7460 12112 7488
rect 12222 7463 12280 7469
rect 12222 7460 12234 7463
rect 12084 7432 12234 7460
rect 8794 7429 8806 7432
rect 8748 7423 8806 7429
rect 12222 7429 12234 7432
rect 12268 7429 12280 7463
rect 13372 7460 13400 7491
rect 13722 7488 13728 7540
rect 13780 7488 13786 7540
rect 13814 7488 13820 7540
rect 13872 7488 13878 7540
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 13832 7460 13860 7488
rect 13372 7432 13860 7460
rect 12222 7423 12280 7429
rect 4430 7352 4436 7404
rect 4488 7352 4494 7404
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 5718 7392 5724 7404
rect 5675 7364 5724 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 3145 7327 3203 7333
rect 3145 7324 3157 7327
rect 2746 7296 3157 7324
rect 3145 7293 3157 7296
rect 3191 7293 3203 7327
rect 3145 7287 3203 7293
rect 3160 7188 3188 7287
rect 3418 7284 3424 7336
rect 3476 7284 3482 7336
rect 4448 7324 4476 7352
rect 5000 7324 5028 7355
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 8481 7395 8539 7401
rect 8481 7361 8493 7395
rect 8527 7392 8539 7395
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 8527 7364 9965 7392
rect 8527 7361 8539 7364
rect 8481 7355 8539 7361
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10220 7395 10278 7401
rect 10220 7361 10232 7395
rect 10266 7392 10278 7395
rect 11054 7392 11060 7404
rect 10266 7364 11060 7392
rect 10266 7361 10278 7364
rect 10220 7355 10278 7361
rect 4448 7296 5028 7324
rect 5902 7284 5908 7336
rect 5960 7284 5966 7336
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7324 7711 7327
rect 7699 7296 8524 7324
rect 7699 7293 7711 7296
rect 7653 7287 7711 7293
rect 4522 7216 4528 7268
rect 4580 7216 4586 7268
rect 4540 7188 4568 7216
rect 8496 7200 8524 7296
rect 3160 7160 4568 7188
rect 5258 7148 5264 7200
rect 5316 7148 5322 7200
rect 8478 7148 8484 7200
rect 8536 7148 8542 7200
rect 9858 7148 9864 7200
rect 9916 7148 9922 7200
rect 9968 7188 9996 7355
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12066 7392 12072 7404
rect 12023 7364 12072 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 13630 7352 13636 7404
rect 13688 7392 13694 7404
rect 14108 7392 14136 7488
rect 15102 7420 15108 7472
rect 15160 7420 15166 7472
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 13688 7364 14044 7392
rect 14108 7364 14197 7392
rect 13688 7352 13694 7364
rect 14016 7324 14044 7364
rect 14185 7361 14197 7364
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7392 15071 7395
rect 15120 7392 15148 7420
rect 15746 7392 15752 7404
rect 15059 7364 15752 7392
rect 15059 7361 15071 7364
rect 15013 7355 15071 7361
rect 15028 7324 15056 7355
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 14016 7296 15056 7324
rect 11256 7228 12020 7256
rect 11256 7188 11284 7228
rect 11992 7200 12020 7228
rect 9968 7160 11284 7188
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 11422 7188 11428 7200
rect 11379 7160 11428 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 11974 7148 11980 7200
rect 12032 7148 12038 7200
rect 13998 7148 14004 7200
rect 14056 7148 14062 7200
rect 15105 7191 15163 7197
rect 15105 7157 15117 7191
rect 15151 7188 15163 7191
rect 15378 7188 15384 7200
rect 15151 7160 15384 7188
rect 15151 7157 15163 7160
rect 15105 7151 15163 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 1104 7098 16652 7120
rect 1104 7046 2893 7098
rect 2945 7046 2957 7098
rect 3009 7046 3021 7098
rect 3073 7046 3085 7098
rect 3137 7046 3149 7098
rect 3201 7046 6780 7098
rect 6832 7046 6844 7098
rect 6896 7046 6908 7098
rect 6960 7046 6972 7098
rect 7024 7046 7036 7098
rect 7088 7046 10667 7098
rect 10719 7046 10731 7098
rect 10783 7046 10795 7098
rect 10847 7046 10859 7098
rect 10911 7046 10923 7098
rect 10975 7046 14554 7098
rect 14606 7046 14618 7098
rect 14670 7046 14682 7098
rect 14734 7046 14746 7098
rect 14798 7046 14810 7098
rect 14862 7046 16652 7098
rect 1104 7024 16652 7046
rect 1670 6944 1676 6996
rect 1728 6944 1734 6996
rect 2590 6984 2596 6996
rect 2516 6956 2596 6984
rect 2516 6857 2544 6956
rect 2590 6944 2596 6956
rect 2648 6944 2654 6996
rect 2774 6984 2780 6996
rect 2746 6944 2780 6984
rect 2832 6944 2838 6996
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3476 6956 3893 6984
rect 3476 6944 3482 6956
rect 3881 6953 3893 6956
rect 3927 6953 3939 6987
rect 3881 6947 3939 6953
rect 11054 6944 11060 6996
rect 11112 6944 11118 6996
rect 13998 6944 14004 6996
rect 14056 6984 14062 6996
rect 14350 6987 14408 6993
rect 14350 6984 14362 6987
rect 14056 6956 14362 6984
rect 14056 6944 14062 6956
rect 14350 6953 14362 6956
rect 14396 6953 14408 6987
rect 14350 6947 14408 6953
rect 2501 6851 2559 6857
rect 2501 6848 2513 6851
rect 2240 6820 2513 6848
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 1872 6644 1900 6743
rect 2240 6712 2268 6820
rect 2501 6817 2513 6820
rect 2547 6817 2559 6851
rect 2746 6848 2774 6944
rect 5350 6876 5356 6928
rect 5408 6916 5414 6928
rect 5902 6916 5908 6928
rect 5408 6888 5908 6916
rect 5408 6876 5414 6888
rect 5902 6876 5908 6888
rect 5960 6916 5966 6928
rect 5960 6888 6224 6916
rect 5960 6876 5966 6888
rect 3418 6848 3424 6860
rect 2501 6811 2559 6817
rect 2608 6820 2774 6848
rect 3068 6820 3424 6848
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 2608 6780 2636 6820
rect 2363 6752 2636 6780
rect 2777 6783 2835 6789
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2777 6749 2789 6783
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 2590 6712 2596 6724
rect 2240 6684 2596 6712
rect 2590 6672 2596 6684
rect 2648 6672 2654 6724
rect 2792 6712 2820 6743
rect 2866 6740 2872 6792
rect 2924 6780 2930 6792
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2924 6752 2973 6780
rect 2924 6740 2930 6752
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 3068 6712 3096 6820
rect 3418 6808 3424 6820
rect 3476 6848 3482 6860
rect 5166 6848 5172 6860
rect 3476 6820 5172 6848
rect 3476 6808 3482 6820
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6780 4123 6783
rect 5258 6780 5264 6792
rect 4111 6752 5264 6780
rect 4111 6749 4123 6752
rect 4065 6743 4123 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 6196 6780 6224 6888
rect 11238 6876 11244 6928
rect 11296 6916 11302 6928
rect 11882 6916 11888 6928
rect 11296 6888 11888 6916
rect 11296 6876 11302 6888
rect 11882 6876 11888 6888
rect 11940 6916 11946 6928
rect 12158 6916 12164 6928
rect 11940 6888 12164 6916
rect 11940 6876 11946 6888
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 7374 6808 7380 6860
rect 7432 6808 7438 6860
rect 7469 6851 7527 6857
rect 7469 6817 7481 6851
rect 7515 6848 7527 6851
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 7515 6820 9505 6848
rect 7515 6817 7527 6820
rect 7469 6811 7527 6817
rect 9493 6817 9505 6820
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 10612 6820 11560 6848
rect 7484 6780 7512 6811
rect 6196 6752 7512 6780
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9858 6780 9864 6792
rect 9447 6752 9864 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 2792 6684 3096 6712
rect 5905 6715 5963 6721
rect 5905 6681 5917 6715
rect 5951 6712 5963 6715
rect 6546 6712 6552 6724
rect 5951 6684 6552 6712
rect 5951 6681 5963 6684
rect 5905 6675 5963 6681
rect 6546 6672 6552 6684
rect 6604 6712 6610 6724
rect 10612 6712 10640 6820
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 11238 6780 11244 6792
rect 10919 6752 11244 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 6604 6684 10640 6712
rect 10689 6715 10747 6721
rect 6604 6672 6610 6684
rect 10689 6681 10701 6715
rect 10735 6681 10747 6715
rect 10689 6675 10747 6681
rect 10781 6715 10839 6721
rect 10781 6681 10793 6715
rect 10827 6712 10839 6715
rect 11422 6712 11428 6724
rect 10827 6684 11428 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 1949 6647 2007 6653
rect 1949 6644 1961 6647
rect 1872 6616 1961 6644
rect 1949 6613 1961 6616
rect 1995 6613 2007 6647
rect 1949 6607 2007 6613
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 3145 6647 3203 6653
rect 3145 6644 3157 6647
rect 2455 6616 3157 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 3145 6613 3157 6616
rect 3191 6613 3203 6647
rect 3145 6607 3203 6613
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 5997 6647 6055 6653
rect 5997 6644 6009 6647
rect 4580 6616 6009 6644
rect 4580 6604 4586 6616
rect 5997 6613 6009 6616
rect 6043 6644 6055 6647
rect 6362 6644 6368 6656
rect 6043 6616 6368 6644
rect 6043 6613 6055 6616
rect 5997 6607 6055 6613
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 6914 6604 6920 6656
rect 6972 6604 6978 6656
rect 7282 6604 7288 6656
rect 7340 6604 7346 6656
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 7616 6616 8953 6644
rect 7616 6604 7622 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 9306 6604 9312 6656
rect 9364 6604 9370 6656
rect 10704 6644 10732 6675
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 11532 6712 11560 6820
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 12342 6848 12348 6860
rect 12032 6820 12348 6848
rect 12032 6808 12038 6820
rect 12342 6808 12348 6820
rect 12400 6848 12406 6860
rect 13906 6848 13912 6860
rect 12400 6820 13912 6848
rect 12400 6808 12406 6820
rect 13906 6808 13912 6820
rect 13964 6848 13970 6860
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13964 6820 14105 6848
rect 13964 6808 13970 6820
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 14093 6811 14151 6817
rect 13725 6715 13783 6721
rect 13725 6712 13737 6715
rect 11532 6684 13737 6712
rect 13725 6681 13737 6684
rect 13771 6712 13783 6715
rect 14274 6712 14280 6724
rect 13771 6684 14280 6712
rect 13771 6681 13783 6684
rect 13725 6675 13783 6681
rect 14274 6672 14280 6684
rect 14332 6672 14338 6724
rect 15378 6672 15384 6724
rect 15436 6672 15442 6724
rect 11146 6644 11152 6656
rect 10704 6616 11152 6644
rect 11146 6604 11152 6616
rect 11204 6644 11210 6656
rect 11790 6644 11796 6656
rect 11204 6616 11796 6644
rect 11204 6604 11210 6616
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 15838 6604 15844 6656
rect 15896 6604 15902 6656
rect 1104 6554 16811 6576
rect 1104 6502 4836 6554
rect 4888 6502 4900 6554
rect 4952 6502 4964 6554
rect 5016 6502 5028 6554
rect 5080 6502 5092 6554
rect 5144 6502 8723 6554
rect 8775 6502 8787 6554
rect 8839 6502 8851 6554
rect 8903 6502 8915 6554
rect 8967 6502 8979 6554
rect 9031 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 16497 6554
rect 16549 6502 16561 6554
rect 16613 6502 16625 6554
rect 16677 6502 16689 6554
rect 16741 6502 16753 6554
rect 16805 6502 16811 6554
rect 1104 6480 16811 6502
rect 6914 6440 6920 6452
rect 3436 6412 6920 6440
rect 3436 6313 3464 6412
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 7282 6400 7288 6452
rect 7340 6440 7346 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 7340 6412 8125 6440
rect 7340 6400 7346 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 8113 6403 8171 6409
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 14645 6443 14703 6449
rect 12299 6412 12434 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 4522 6372 4528 6384
rect 4264 6344 4528 6372
rect 4264 6313 4292 6344
rect 4522 6332 4528 6344
rect 4580 6332 4586 6384
rect 5258 6332 5264 6384
rect 5316 6332 5322 6384
rect 7098 6332 7104 6384
rect 7156 6332 7162 6384
rect 9490 6332 9496 6384
rect 9548 6372 9554 6384
rect 12406 6372 12434 6412
rect 14645 6409 14657 6443
rect 14691 6440 14703 6443
rect 15838 6440 15844 6452
rect 14691 6412 15844 6440
rect 14691 6409 14703 6412
rect 14645 6403 14703 6409
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 12590 6375 12648 6381
rect 12590 6372 12602 6375
rect 9548 6344 12296 6372
rect 12406 6344 12602 6372
rect 9548 6332 9554 6344
rect 12268 6316 12296 6344
rect 12590 6341 12602 6344
rect 12636 6341 12648 6375
rect 12590 6335 12648 6341
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 11330 6264 11336 6316
rect 11388 6304 11394 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11388 6276 11713 6304
rect 11388 6264 11394 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11790 6264 11796 6316
rect 11848 6304 11854 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11848 6276 11897 6304
rect 11848 6264 11854 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6304 12127 6307
rect 12158 6304 12164 6316
rect 12115 6276 12164 6304
rect 12115 6273 12127 6276
rect 12069 6267 12127 6273
rect 4522 6196 4528 6248
rect 4580 6196 4586 6248
rect 5718 6196 5724 6248
rect 5776 6196 5782 6248
rect 6638 6196 6644 6248
rect 6696 6196 6702 6248
rect 5736 6168 5764 6196
rect 5997 6171 6055 6177
rect 5997 6168 6009 6171
rect 5736 6140 6009 6168
rect 5997 6137 6009 6140
rect 6043 6137 6055 6171
rect 5997 6131 6055 6137
rect 3234 6060 3240 6112
rect 3292 6060 3298 6112
rect 8662 6060 8668 6112
rect 8720 6060 8726 6112
rect 11992 6100 12020 6267
rect 12158 6264 12164 6276
rect 12216 6264 12222 6316
rect 12250 6264 12256 6316
rect 12308 6264 12314 6316
rect 12342 6196 12348 6248
rect 12400 6196 12406 6248
rect 14737 6239 14795 6245
rect 14737 6205 14749 6239
rect 14783 6205 14795 6239
rect 14737 6199 14795 6205
rect 13725 6171 13783 6177
rect 13725 6137 13737 6171
rect 13771 6168 13783 6171
rect 14752 6168 14780 6199
rect 14918 6196 14924 6248
rect 14976 6196 14982 6248
rect 13771 6140 14780 6168
rect 13771 6137 13783 6140
rect 13725 6131 13783 6137
rect 13740 6100 13768 6131
rect 11992 6072 13768 6100
rect 14274 6060 14280 6112
rect 14332 6060 14338 6112
rect 1104 6010 16652 6032
rect 1104 5958 2893 6010
rect 2945 5958 2957 6010
rect 3009 5958 3021 6010
rect 3073 5958 3085 6010
rect 3137 5958 3149 6010
rect 3201 5958 6780 6010
rect 6832 5958 6844 6010
rect 6896 5958 6908 6010
rect 6960 5958 6972 6010
rect 7024 5958 7036 6010
rect 7088 5958 10667 6010
rect 10719 5958 10731 6010
rect 10783 5958 10795 6010
rect 10847 5958 10859 6010
rect 10911 5958 10923 6010
rect 10975 5958 14554 6010
rect 14606 5958 14618 6010
rect 14670 5958 14682 6010
rect 14734 5958 14746 6010
rect 14798 5958 14810 6010
rect 14862 5958 16652 6010
rect 1104 5936 16652 5958
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3418 5896 3424 5908
rect 3016 5868 3424 5896
rect 3016 5856 3022 5868
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 4522 5856 4528 5908
rect 4580 5896 4586 5908
rect 4801 5899 4859 5905
rect 4801 5896 4813 5899
rect 4580 5868 4813 5896
rect 4580 5856 4586 5868
rect 4801 5865 4813 5868
rect 4847 5865 4859 5899
rect 4801 5859 4859 5865
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5316 5868 5365 5896
rect 5316 5856 5322 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 6181 5899 6239 5905
rect 6181 5865 6193 5899
rect 6227 5896 6239 5899
rect 6638 5896 6644 5908
rect 6227 5868 6644 5896
rect 6227 5865 6239 5868
rect 6181 5859 6239 5865
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5896 6883 5899
rect 7098 5896 7104 5908
rect 6871 5868 7104 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 8662 5856 8668 5908
rect 8720 5856 8726 5908
rect 8846 5856 8852 5908
rect 8904 5896 8910 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8904 5868 9137 5896
rect 8904 5856 8910 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 9306 5856 9312 5908
rect 9364 5856 9370 5908
rect 10244 5868 12112 5896
rect 6454 5788 6460 5840
rect 6512 5828 6518 5840
rect 6512 5800 7052 5828
rect 6512 5788 6518 5800
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 3326 5760 3332 5772
rect 2731 5732 3332 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 5442 5760 5448 5772
rect 5276 5732 5448 5760
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2832 5664 2881 5692
rect 2832 5652 2838 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 3881 5695 3939 5701
rect 3881 5661 3893 5695
rect 3927 5692 3939 5695
rect 4430 5692 4436 5704
rect 3927 5664 4436 5692
rect 3927 5661 3939 5664
rect 3881 5655 3939 5661
rect 2884 5624 2912 5655
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5692 5043 5695
rect 5166 5692 5172 5704
rect 5031 5664 5172 5692
rect 5031 5661 5043 5664
rect 4985 5655 5043 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5276 5701 5304 5732
rect 5442 5720 5448 5732
rect 5500 5760 5506 5772
rect 7024 5769 7052 5800
rect 7009 5763 7067 5769
rect 5500 5732 6776 5760
rect 5500 5720 5506 5732
rect 6748 5701 6776 5732
rect 7009 5729 7021 5763
rect 7055 5729 7067 5763
rect 7009 5723 7067 5729
rect 7285 5763 7343 5769
rect 7285 5729 7297 5763
rect 7331 5760 7343 5763
rect 8680 5760 8708 5856
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 9324 5828 9352 5856
rect 8803 5800 9352 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 7331 5732 8708 5760
rect 7331 5729 7343 5732
rect 7285 5723 7343 5729
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9548 5732 9689 5760
rect 9548 5720 9554 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5760 10195 5763
rect 10244 5760 10272 5868
rect 12084 5840 12112 5868
rect 12250 5856 12256 5908
rect 12308 5896 12314 5908
rect 12308 5868 12572 5896
rect 12308 5856 12314 5868
rect 12066 5788 12072 5840
rect 12124 5788 12130 5840
rect 10183 5732 10272 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 11422 5720 11428 5772
rect 11480 5760 11486 5772
rect 12544 5769 12572 5868
rect 14274 5856 14280 5908
rect 14332 5856 14338 5908
rect 16114 5856 16120 5908
rect 16172 5856 16178 5908
rect 12437 5763 12495 5769
rect 12437 5760 12449 5763
rect 11480 5732 12449 5760
rect 11480 5720 11486 5732
rect 12437 5729 12449 5732
rect 12483 5729 12495 5763
rect 12437 5723 12495 5729
rect 12529 5763 12587 5769
rect 12529 5729 12541 5763
rect 12575 5729 12587 5763
rect 12529 5723 12587 5729
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5661 6791 5695
rect 6733 5655 6791 5661
rect 4062 5624 4068 5636
rect 2884 5596 4068 5624
rect 4062 5584 4068 5596
rect 4120 5584 4126 5636
rect 4448 5624 4476 5652
rect 5276 5624 5304 5655
rect 4448 5596 5304 5624
rect 6380 5624 6408 5655
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 12805 5695 12863 5701
rect 12805 5692 12817 5695
rect 12676 5664 12817 5692
rect 12676 5652 12682 5664
rect 12805 5661 12817 5664
rect 12851 5692 12863 5695
rect 13630 5692 13636 5704
rect 12851 5664 13636 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 14292 5692 14320 5856
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14292 5664 14565 5692
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5692 16359 5695
rect 16347 5664 16988 5692
rect 16347 5661 16359 5664
rect 16301 5655 16359 5661
rect 16960 5636 16988 5664
rect 7558 5624 7564 5636
rect 6380 5596 7564 5624
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 8294 5584 8300 5636
rect 8352 5584 8358 5636
rect 9493 5627 9551 5633
rect 9493 5593 9505 5627
rect 9539 5624 9551 5627
rect 9539 5596 10364 5624
rect 9539 5593 9551 5596
rect 9493 5587 9551 5593
rect 3050 5516 3056 5568
rect 3108 5516 3114 5568
rect 3970 5516 3976 5568
rect 4028 5516 4034 5568
rect 9582 5516 9588 5568
rect 9640 5516 9646 5568
rect 10336 5556 10364 5596
rect 10410 5584 10416 5636
rect 10468 5584 10474 5636
rect 12897 5627 12955 5633
rect 12897 5624 12909 5627
rect 11638 5596 12909 5624
rect 12897 5593 12909 5596
rect 12943 5593 12955 5627
rect 12897 5587 12955 5593
rect 16942 5584 16948 5636
rect 17000 5584 17006 5636
rect 11885 5559 11943 5565
rect 11885 5556 11897 5559
rect 10336 5528 11897 5556
rect 11885 5525 11897 5528
rect 11931 5525 11943 5559
rect 11885 5519 11943 5525
rect 11974 5516 11980 5568
rect 12032 5516 12038 5568
rect 12342 5516 12348 5568
rect 12400 5516 12406 5568
rect 14366 5516 14372 5568
rect 14424 5516 14430 5568
rect 1104 5466 16811 5488
rect 1104 5414 4836 5466
rect 4888 5414 4900 5466
rect 4952 5414 4964 5466
rect 5016 5414 5028 5466
rect 5080 5414 5092 5466
rect 5144 5414 8723 5466
rect 8775 5414 8787 5466
rect 8839 5414 8851 5466
rect 8903 5414 8915 5466
rect 8967 5414 8979 5466
rect 9031 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 16497 5466
rect 16549 5414 16561 5466
rect 16613 5414 16625 5466
rect 16677 5414 16689 5466
rect 16741 5414 16753 5466
rect 16805 5414 16811 5466
rect 1104 5392 16811 5414
rect 1857 5355 1915 5361
rect 1857 5321 1869 5355
rect 1903 5321 1915 5355
rect 1857 5315 1915 5321
rect 2317 5355 2375 5361
rect 2317 5321 2329 5355
rect 2363 5352 2375 5355
rect 3050 5352 3056 5364
rect 2363 5324 3056 5352
rect 2363 5321 2375 5324
rect 2317 5315 2375 5321
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 1872 5216 1900 5315
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8294 5352 8300 5364
rect 7975 5324 8300 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 9582 5312 9588 5364
rect 9640 5352 9646 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9640 5324 10057 5352
rect 9640 5312 9646 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10045 5315 10103 5321
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 10468 5324 10517 5352
rect 10468 5312 10474 5324
rect 10505 5321 10517 5324
rect 10551 5321 10563 5355
rect 10505 5315 10563 5321
rect 11974 5312 11980 5364
rect 12032 5312 12038 5364
rect 12161 5355 12219 5361
rect 12161 5321 12173 5355
rect 12207 5352 12219 5355
rect 12207 5324 12434 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 2225 5287 2283 5293
rect 2225 5253 2237 5287
rect 2271 5284 2283 5287
rect 2498 5284 2504 5296
rect 2271 5256 2504 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 2498 5244 2504 5256
rect 2556 5244 2562 5296
rect 2961 5287 3019 5293
rect 2961 5253 2973 5287
rect 3007 5284 3019 5287
rect 3234 5284 3240 5296
rect 3007 5256 3240 5284
rect 3007 5253 3019 5256
rect 2961 5247 3019 5253
rect 3234 5244 3240 5256
rect 3292 5244 3298 5296
rect 3970 5244 3976 5296
rect 4028 5244 4034 5296
rect 9490 5284 9496 5296
rect 8680 5256 9496 5284
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 1811 5188 1900 5216
rect 2424 5188 2697 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 2424 5160 2452 5188
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 4706 5176 4712 5228
rect 4764 5216 4770 5228
rect 8680 5225 8708 5256
rect 9490 5244 9496 5256
rect 9548 5244 9554 5296
rect 11992 5284 12020 5312
rect 10704 5256 12020 5284
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 4764 5188 5457 5216
rect 4764 5176 4770 5188
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 5445 5179 5503 5185
rect 7392 5188 7849 5216
rect 2406 5108 2412 5160
rect 2464 5108 2470 5160
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 2590 5148 2596 5160
rect 2547 5120 2596 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 7392 5024 7420 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 8932 5219 8990 5225
rect 8932 5185 8944 5219
rect 8978 5216 8990 5219
rect 9766 5216 9772 5228
rect 8978 5188 9772 5216
rect 8978 5185 8990 5188
rect 8932 5179 8990 5185
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 10704 5225 10732 5256
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 12406 5284 12434 5324
rect 12498 5287 12556 5293
rect 12498 5284 12510 5287
rect 12124 5256 12296 5284
rect 12406 5256 12510 5284
rect 12124 5244 12130 5256
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 11606 5176 11612 5228
rect 11664 5176 11670 5228
rect 11790 5176 11796 5228
rect 11848 5176 11854 5228
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12158 5216 12164 5228
rect 12023 5188 12164 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 1670 5012 1676 5024
rect 1627 4984 1676 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 4433 5015 4491 5021
rect 4433 5012 4445 5015
rect 4212 4984 4445 5012
rect 4212 4972 4218 4984
rect 4433 4981 4445 4984
rect 4479 4981 4491 5015
rect 4433 4975 4491 4981
rect 5258 4972 5264 5024
rect 5316 4972 5322 5024
rect 7374 4972 7380 5024
rect 7432 4972 7438 5024
rect 11900 5012 11928 5179
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12268 5225 12296 5256
rect 12498 5253 12510 5256
rect 12544 5253 12556 5287
rect 12498 5247 12556 5253
rect 14366 5244 14372 5296
rect 14424 5284 14430 5296
rect 14461 5287 14519 5293
rect 14461 5284 14473 5287
rect 14424 5256 14473 5284
rect 14424 5244 14430 5256
rect 14461 5253 14473 5256
rect 14507 5253 14519 5287
rect 16117 5287 16175 5293
rect 16117 5284 16129 5287
rect 15686 5256 16129 5284
rect 14461 5247 14519 5253
rect 16117 5253 16129 5256
rect 16163 5253 16175 5287
rect 16117 5247 16175 5253
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 13906 5216 13912 5228
rect 12299 5188 13912 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 13906 5176 13912 5188
rect 13964 5216 13970 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 13964 5188 14197 5216
rect 13964 5176 13970 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 15746 5176 15752 5228
rect 15804 5216 15810 5228
rect 16025 5219 16083 5225
rect 16025 5216 16037 5219
rect 15804 5188 16037 5216
rect 15804 5176 15810 5188
rect 16025 5185 16037 5188
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 13630 5012 13636 5024
rect 11900 4984 13636 5012
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 15930 4972 15936 5024
rect 15988 4972 15994 5024
rect 1104 4922 16652 4944
rect 1104 4870 2893 4922
rect 2945 4870 2957 4922
rect 3009 4870 3021 4922
rect 3073 4870 3085 4922
rect 3137 4870 3149 4922
rect 3201 4870 6780 4922
rect 6832 4870 6844 4922
rect 6896 4870 6908 4922
rect 6960 4870 6972 4922
rect 7024 4870 7036 4922
rect 7088 4870 10667 4922
rect 10719 4870 10731 4922
rect 10783 4870 10795 4922
rect 10847 4870 10859 4922
rect 10911 4870 10923 4922
rect 10975 4870 14554 4922
rect 14606 4870 14618 4922
rect 14670 4870 14682 4922
rect 14734 4870 14746 4922
rect 14798 4870 14810 4922
rect 14862 4870 16652 4922
rect 1104 4848 16652 4870
rect 4706 4768 4712 4820
rect 4764 4768 4770 4820
rect 5258 4768 5264 4820
rect 5316 4768 5322 4820
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 7374 4808 7380 4820
rect 5500 4780 7380 4808
rect 5500 4768 5506 4780
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 9766 4768 9772 4820
rect 9824 4768 9830 4820
rect 13630 4768 13636 4820
rect 13688 4768 13694 4820
rect 15930 4768 15936 4820
rect 15988 4768 15994 4820
rect 2498 4700 2504 4752
rect 2556 4740 2562 4752
rect 2777 4743 2835 4749
rect 2777 4740 2789 4743
rect 2556 4712 2789 4740
rect 2556 4700 2562 4712
rect 2777 4709 2789 4712
rect 2823 4740 2835 4743
rect 5276 4740 5304 4768
rect 2823 4712 3464 4740
rect 5276 4712 5580 4740
rect 2823 4709 2835 4712
rect 2777 4703 2835 4709
rect 1670 4613 1676 4616
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4573 1455 4607
rect 1664 4604 1676 4613
rect 1631 4576 1676 4604
rect 1397 4567 1455 4573
rect 1664 4567 1676 4576
rect 1412 4536 1440 4567
rect 1670 4564 1676 4567
rect 1728 4564 1734 4616
rect 2406 4564 2412 4616
rect 2464 4564 2470 4616
rect 2424 4536 2452 4564
rect 1412 4508 2452 4536
rect 3436 4536 3464 4712
rect 5350 4632 5356 4684
rect 5408 4632 5414 4684
rect 5552 4672 5580 4712
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 5552 4644 5825 4672
rect 5813 4641 5825 4644
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4430 4604 4436 4616
rect 4387 4576 4436 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4604 5135 4607
rect 5166 4604 5172 4616
rect 5123 4576 5172 4604
rect 5123 4573 5135 4576
rect 5077 4567 5135 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 7392 4613 7420 4768
rect 13648 4672 13676 4768
rect 13814 4700 13820 4752
rect 13872 4740 13878 4752
rect 13872 4712 14780 4740
rect 13872 4700 13878 4712
rect 14752 4681 14780 4712
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 9416 4644 11836 4672
rect 13648 4644 14565 4672
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 7423 4576 7665 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 3436 4508 5212 4536
rect 3786 4428 3792 4480
rect 3844 4428 3850 4480
rect 4430 4428 4436 4480
rect 4488 4428 4494 4480
rect 5184 4477 5212 4508
rect 5169 4471 5227 4477
rect 5169 4437 5181 4471
rect 5215 4437 5227 4471
rect 5552 4468 5580 4567
rect 9214 4564 9220 4616
rect 9272 4564 9278 4616
rect 9416 4613 9444 4644
rect 11808 4616 11836 4644
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 14918 4672 14924 4684
rect 14783 4644 14924 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 14918 4632 14924 4644
rect 14976 4632 14982 4684
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 7469 4539 7527 4545
rect 7469 4536 7481 4539
rect 7038 4508 7481 4536
rect 7469 4505 7481 4508
rect 7515 4505 7527 4539
rect 7469 4499 7527 4505
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4505 9551 4539
rect 9600 4536 9628 4567
rect 10318 4564 10324 4616
rect 10376 4564 10382 4616
rect 11790 4564 11796 4616
rect 11848 4564 11854 4616
rect 12158 4564 12164 4616
rect 12216 4564 12222 4616
rect 13909 4607 13967 4613
rect 13909 4573 13921 4607
rect 13955 4604 13967 4607
rect 14461 4607 14519 4613
rect 13955 4576 14136 4604
rect 13955 4573 13967 4576
rect 13909 4567 13967 4573
rect 12176 4536 12204 4564
rect 9600 4508 12204 4536
rect 9493 4499 9551 4505
rect 6454 4468 6460 4480
rect 5552 4440 6460 4468
rect 5169 4431 5227 4437
rect 6454 4428 6460 4440
rect 6512 4428 6518 4480
rect 7282 4428 7288 4480
rect 7340 4428 7346 4480
rect 7742 4428 7748 4480
rect 7800 4428 7806 4480
rect 9508 4468 9536 4499
rect 9582 4468 9588 4480
rect 9508 4440 9588 4468
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 10134 4428 10140 4480
rect 10192 4428 10198 4480
rect 13725 4471 13783 4477
rect 13725 4437 13737 4471
rect 13771 4468 13783 4471
rect 13998 4468 14004 4480
rect 13771 4440 14004 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 14108 4477 14136 4576
rect 14461 4573 14473 4607
rect 14507 4604 14519 4607
rect 15948 4604 15976 4768
rect 14507 4576 15976 4604
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 14093 4471 14151 4477
rect 14093 4437 14105 4471
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 1104 4378 16811 4400
rect 1104 4326 4836 4378
rect 4888 4326 4900 4378
rect 4952 4326 4964 4378
rect 5016 4326 5028 4378
rect 5080 4326 5092 4378
rect 5144 4326 8723 4378
rect 8775 4326 8787 4378
rect 8839 4326 8851 4378
rect 8903 4326 8915 4378
rect 8967 4326 8979 4378
rect 9031 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 16497 4378
rect 16549 4326 16561 4378
rect 16613 4326 16625 4378
rect 16677 4326 16689 4378
rect 16741 4326 16753 4378
rect 16805 4326 16811 4378
rect 1104 4304 16811 4326
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 5629 4267 5687 4273
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 5675 4236 8493 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8481 4227 8539 4233
rect 13081 4267 13139 4273
rect 13081 4233 13093 4267
rect 13127 4264 13139 4267
rect 15473 4267 15531 4273
rect 15473 4264 15485 4267
rect 13127 4236 15485 4264
rect 13127 4233 13139 4236
rect 13081 4227 13139 4233
rect 15473 4233 15485 4236
rect 15519 4233 15531 4267
rect 15473 4227 15531 4233
rect 934 4156 940 4208
rect 992 4196 998 4208
rect 1489 4199 1547 4205
rect 1489 4196 1501 4199
rect 992 4168 1501 4196
rect 992 4156 998 4168
rect 1489 4165 1501 4168
rect 1535 4165 1547 4199
rect 1489 4159 1547 4165
rect 3697 4199 3755 4205
rect 3697 4165 3709 4199
rect 3743 4196 3755 4199
rect 3786 4196 3792 4208
rect 3743 4168 3792 4196
rect 3743 4165 3755 4168
rect 3697 4159 3755 4165
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 4430 4156 4436 4208
rect 4488 4156 4494 4208
rect 7742 4156 7748 4208
rect 7800 4156 7806 4208
rect 9861 4199 9919 4205
rect 9861 4165 9873 4199
rect 9907 4196 9919 4199
rect 10134 4196 10140 4208
rect 9907 4168 10140 4196
rect 9907 4165 9919 4168
rect 9861 4159 9919 4165
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 13906 4196 13912 4208
rect 11086 4168 11652 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 2774 4128 2780 4140
rect 1719 4100 2780 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 6454 4128 6460 4140
rect 5460 4100 6460 4128
rect 2406 4020 2412 4072
rect 2464 4060 2470 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 2464 4032 3433 4060
rect 2464 4020 2470 4032
rect 3421 4029 3433 4032
rect 3467 4060 3479 4063
rect 5460 4060 5488 4100
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 6638 4088 6644 4140
rect 6696 4088 6702 4140
rect 11514 4088 11520 4140
rect 11572 4088 11578 4140
rect 11624 4137 11652 4168
rect 12176 4168 12388 4196
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 3467 4032 5488 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 5718 4020 5724 4072
rect 5776 4020 5782 4072
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4029 5871 4063
rect 6472 4060 6500 4088
rect 6733 4063 6791 4069
rect 6733 4060 6745 4063
rect 6472 4032 6745 4060
rect 5813 4023 5871 4029
rect 6733 4029 6745 4032
rect 6779 4029 6791 4063
rect 7009 4063 7067 4069
rect 7009 4060 7021 4063
rect 6733 4023 6791 4029
rect 6840 4032 7021 4060
rect 5350 3992 5356 4004
rect 5184 3964 5356 3992
rect 4430 3884 4436 3936
rect 4488 3924 4494 3936
rect 5184 3924 5212 3964
rect 5350 3952 5356 3964
rect 5408 3992 5414 4004
rect 5828 3992 5856 4023
rect 5408 3964 5856 3992
rect 6457 3995 6515 4001
rect 5408 3952 5414 3964
rect 6457 3961 6469 3995
rect 6503 3992 6515 3995
rect 6840 3992 6868 4032
rect 7009 4029 7021 4032
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 9582 4020 9588 4072
rect 9640 4020 9646 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 12176 4060 12204 4168
rect 12360 4140 12388 4168
rect 13740 4168 13912 4196
rect 12250 4088 12256 4140
rect 12308 4088 12314 4140
rect 12342 4088 12348 4140
rect 12400 4088 12406 4140
rect 13740 4137 13768 4168
rect 13906 4156 13912 4168
rect 13964 4156 13970 4208
rect 15226 4168 15700 4196
rect 15672 4137 15700 4168
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 13725 4131 13783 4137
rect 12575 4100 12756 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 11379 4032 12204 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 6503 3964 6868 3992
rect 6503 3961 6515 3964
rect 6457 3955 6515 3961
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 12268 3992 12296 4088
rect 12728 4001 12756 4100
rect 13725 4097 13737 4131
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4097 15623 4131
rect 15565 4091 15623 4097
rect 15657 4131 15715 4137
rect 15657 4097 15669 4131
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 13170 4020 13176 4072
rect 13228 4020 13234 4072
rect 13357 4063 13415 4069
rect 13357 4029 13369 4063
rect 13403 4060 13415 4063
rect 13403 4032 13768 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 12713 3995 12771 4001
rect 11112 3964 12664 3992
rect 11112 3952 11118 3964
rect 4488 3896 5212 3924
rect 4488 3884 4494 3896
rect 5258 3884 5264 3936
rect 5316 3884 5322 3936
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 12308 3896 12357 3924
rect 12308 3884 12314 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12636 3924 12664 3964
rect 12713 3961 12725 3995
rect 12759 3961 12771 3995
rect 12713 3955 12771 3961
rect 13372 3924 13400 4023
rect 13740 4004 13768 4032
rect 13998 4020 14004 4072
rect 14056 4020 14062 4072
rect 15580 4060 15608 4091
rect 15746 4060 15752 4072
rect 15580 4032 15752 4060
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 13722 3952 13728 4004
rect 13780 3952 13786 4004
rect 12636 3896 13400 3924
rect 12345 3887 12403 3893
rect 1104 3834 16652 3856
rect 1104 3782 2893 3834
rect 2945 3782 2957 3834
rect 3009 3782 3021 3834
rect 3073 3782 3085 3834
rect 3137 3782 3149 3834
rect 3201 3782 6780 3834
rect 6832 3782 6844 3834
rect 6896 3782 6908 3834
rect 6960 3782 6972 3834
rect 7024 3782 7036 3834
rect 7088 3782 10667 3834
rect 10719 3782 10731 3834
rect 10783 3782 10795 3834
rect 10847 3782 10859 3834
rect 10911 3782 10923 3834
rect 10975 3782 14554 3834
rect 14606 3782 14618 3834
rect 14670 3782 14682 3834
rect 14734 3782 14746 3834
rect 14798 3782 14810 3834
rect 14862 3782 16652 3834
rect 1104 3760 16652 3782
rect 3789 3723 3847 3729
rect 3789 3689 3801 3723
rect 3835 3720 3847 3723
rect 3970 3720 3976 3732
rect 3835 3692 3976 3720
rect 3835 3689 3847 3692
rect 3789 3683 3847 3689
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 6638 3680 6644 3732
rect 6696 3720 6702 3732
rect 7009 3723 7067 3729
rect 7009 3720 7021 3723
rect 6696 3692 7021 3720
rect 6696 3680 6702 3692
rect 7009 3689 7021 3692
rect 7055 3689 7067 3723
rect 7009 3683 7067 3689
rect 10318 3680 10324 3732
rect 10376 3680 10382 3732
rect 11054 3680 11060 3732
rect 11112 3680 11118 3732
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 12526 3720 12532 3732
rect 11572 3692 12532 3720
rect 11572 3680 11578 3692
rect 12526 3680 12532 3692
rect 12584 3720 12590 3732
rect 12584 3692 13768 3720
rect 12584 3680 12590 3692
rect 4430 3544 4436 3596
rect 4488 3584 4494 3596
rect 7561 3587 7619 3593
rect 7561 3584 7573 3587
rect 4488 3556 7573 3584
rect 4488 3544 4494 3556
rect 7561 3553 7573 3556
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3584 11023 3587
rect 11072 3584 11100 3680
rect 11011 3556 11100 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11882 3544 11888 3596
rect 11940 3544 11946 3596
rect 12161 3587 12219 3593
rect 12161 3553 12173 3587
rect 12207 3584 12219 3587
rect 12250 3584 12256 3596
rect 12207 3556 12256 3584
rect 12207 3553 12219 3556
rect 12161 3547 12219 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 2958 3476 2964 3528
rect 3016 3476 3022 3528
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4706 3476 4712 3528
rect 4764 3516 4770 3528
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4764 3488 4905 3516
rect 4764 3476 4770 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 5166 3476 5172 3528
rect 5224 3476 5230 3528
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 5276 3448 5304 3479
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 13740 3525 13768 3692
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 13964 3692 14657 3720
rect 13964 3680 13970 3692
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 14645 3683 14703 3689
rect 14182 3612 14188 3664
rect 14240 3652 14246 3664
rect 14277 3655 14335 3661
rect 14277 3652 14289 3655
rect 14240 3624 14289 3652
rect 14240 3612 14246 3624
rect 14277 3621 14289 3624
rect 14323 3621 14335 3655
rect 14277 3615 14335 3621
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 7340 3488 7389 3516
rect 7340 3476 7346 3488
rect 7377 3485 7389 3488
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3485 14151 3519
rect 14292 3516 14320 3615
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14292 3488 14473 3516
rect 14093 3479 14151 3485
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 8294 3448 8300 3460
rect 4120 3420 8300 3448
rect 4120 3408 4126 3420
rect 8294 3408 8300 3420
rect 8352 3448 8358 3460
rect 8570 3448 8576 3460
rect 8352 3420 8576 3448
rect 8352 3408 8358 3420
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 13817 3451 13875 3457
rect 13817 3448 13829 3451
rect 10704 3420 12434 3448
rect 13386 3420 13829 3448
rect 2774 3340 2780 3392
rect 2832 3340 2838 3392
rect 3786 3340 3792 3392
rect 3844 3380 3850 3392
rect 4249 3383 4307 3389
rect 4249 3380 4261 3383
rect 3844 3352 4261 3380
rect 3844 3340 3850 3352
rect 4249 3349 4261 3352
rect 4295 3349 4307 3383
rect 4249 3343 4307 3349
rect 4706 3340 4712 3392
rect 4764 3340 4770 3392
rect 5442 3340 5448 3392
rect 5500 3340 5506 3392
rect 7466 3340 7472 3392
rect 7524 3340 7530 3392
rect 10704 3389 10732 3420
rect 10689 3383 10747 3389
rect 10689 3349 10701 3383
rect 10735 3349 10747 3383
rect 10689 3343 10747 3349
rect 10778 3340 10784 3392
rect 10836 3340 10842 3392
rect 12406 3380 12434 3420
rect 13817 3417 13829 3420
rect 13863 3417 13875 3451
rect 14108 3448 14136 3479
rect 16114 3448 16120 3460
rect 14108 3420 16120 3448
rect 13817 3411 13875 3417
rect 16114 3408 16120 3420
rect 16172 3408 16178 3460
rect 13633 3383 13691 3389
rect 13633 3380 13645 3383
rect 12406 3352 13645 3380
rect 13633 3349 13645 3352
rect 13679 3349 13691 3383
rect 13633 3343 13691 3349
rect 1104 3290 16811 3312
rect 1104 3238 4836 3290
rect 4888 3238 4900 3290
rect 4952 3238 4964 3290
rect 5016 3238 5028 3290
rect 5080 3238 5092 3290
rect 5144 3238 8723 3290
rect 8775 3238 8787 3290
rect 8839 3238 8851 3290
rect 8903 3238 8915 3290
rect 8967 3238 8979 3290
rect 9031 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 16497 3290
rect 16549 3238 16561 3290
rect 16613 3238 16625 3290
rect 16677 3238 16689 3290
rect 16741 3238 16753 3290
rect 16805 3238 16811 3290
rect 1104 3216 16811 3238
rect 2774 3136 2780 3188
rect 2832 3136 2838 3188
rect 3786 3136 3792 3188
rect 3844 3136 3850 3188
rect 4062 3136 4068 3188
rect 4120 3136 4126 3188
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 5813 3179 5871 3185
rect 5813 3176 5825 3179
rect 5776 3148 5825 3176
rect 5776 3136 5782 3148
rect 5813 3145 5825 3148
rect 5859 3145 5871 3179
rect 5813 3139 5871 3145
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7524 3148 7849 3176
rect 7524 3136 7530 3148
rect 7837 3145 7849 3148
rect 7883 3176 7895 3179
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 7883 3148 8309 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8297 3145 8309 3148
rect 8343 3145 8355 3179
rect 11698 3176 11704 3188
rect 8297 3139 8355 3145
rect 9508 3148 11704 3176
rect 2676 3111 2734 3117
rect 2676 3077 2688 3111
rect 2722 3108 2734 3111
rect 2792 3108 2820 3136
rect 2722 3080 2820 3108
rect 2722 3077 2734 3080
rect 2676 3071 2734 3077
rect 2406 3000 2412 3052
rect 2464 3000 2470 3052
rect 3878 3000 3884 3052
rect 3936 3000 3942 3052
rect 4080 3049 4108 3136
rect 4706 3117 4712 3120
rect 4689 3111 4712 3117
rect 4689 3077 4701 3111
rect 4689 3071 4712 3077
rect 4706 3068 4712 3071
rect 4764 3068 4770 3120
rect 8389 3111 8447 3117
rect 8389 3077 8401 3111
rect 8435 3108 8447 3111
rect 9125 3111 9183 3117
rect 9125 3108 9137 3111
rect 8435 3080 9137 3108
rect 8435 3077 8447 3080
rect 8389 3071 8447 3077
rect 9125 3077 9137 3080
rect 9171 3077 9183 3111
rect 9125 3071 9183 3077
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 6454 3040 6460 3052
rect 4479 3012 6460 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 6724 3043 6782 3049
rect 6724 3009 6736 3043
rect 6770 3040 6782 3043
rect 7098 3040 7104 3052
rect 6770 3012 7104 3040
rect 6770 3009 6782 3012
rect 6724 3003 6782 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8352 3012 8953 3040
rect 8352 3000 8358 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 8478 2932 8484 2984
rect 8536 2932 8542 2984
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 9508 2972 9536 3148
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 13357 3179 13415 3185
rect 13357 3176 13369 3179
rect 13228 3148 13369 3176
rect 13228 3136 13234 3148
rect 13357 3145 13369 3148
rect 13403 3145 13415 3179
rect 13357 3139 13415 3145
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 9640 3080 11928 3108
rect 9640 3068 9646 3080
rect 9784 3049 9812 3080
rect 11900 3052 11928 3080
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 10036 3043 10094 3049
rect 10036 3009 10048 3043
rect 10082 3040 10094 3043
rect 10502 3040 10508 3052
rect 10082 3012 10508 3040
rect 10082 3009 10094 3012
rect 10036 3003 10094 3009
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 11882 3000 11888 3052
rect 11940 3040 11946 3052
rect 12250 3049 12256 3052
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11940 3012 11989 3040
rect 11940 3000 11946 3012
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12244 3003 12256 3049
rect 12250 3000 12256 3003
rect 12308 3000 12314 3052
rect 8803 2944 9536 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 4246 2796 4252 2848
rect 4304 2796 4310 2848
rect 7926 2796 7932 2848
rect 7984 2796 7990 2848
rect 10410 2796 10416 2848
rect 10468 2836 10474 2848
rect 10778 2836 10784 2848
rect 10468 2808 10784 2836
rect 10468 2796 10474 2808
rect 10778 2796 10784 2808
rect 10836 2836 10842 2848
rect 11149 2839 11207 2845
rect 11149 2836 11161 2839
rect 10836 2808 11161 2836
rect 10836 2796 10842 2808
rect 11149 2805 11161 2808
rect 11195 2805 11207 2839
rect 11149 2799 11207 2805
rect 1104 2746 16652 2768
rect 1104 2694 2893 2746
rect 2945 2694 2957 2746
rect 3009 2694 3021 2746
rect 3073 2694 3085 2746
rect 3137 2694 3149 2746
rect 3201 2694 6780 2746
rect 6832 2694 6844 2746
rect 6896 2694 6908 2746
rect 6960 2694 6972 2746
rect 7024 2694 7036 2746
rect 7088 2694 10667 2746
rect 10719 2694 10731 2746
rect 10783 2694 10795 2746
rect 10847 2694 10859 2746
rect 10911 2694 10923 2746
rect 10975 2694 14554 2746
rect 14606 2694 14618 2746
rect 14670 2694 14682 2746
rect 14734 2694 14746 2746
rect 14798 2694 14810 2746
rect 14862 2694 16652 2746
rect 1104 2672 16652 2694
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 2869 2635 2927 2641
rect 2869 2632 2881 2635
rect 2832 2604 2881 2632
rect 2832 2592 2838 2604
rect 2869 2601 2881 2604
rect 2915 2601 2927 2635
rect 2869 2595 2927 2601
rect 3878 2592 3884 2644
rect 3936 2592 3942 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 4893 2635 4951 2641
rect 4893 2632 4905 2635
rect 4764 2604 4905 2632
rect 4764 2592 4770 2604
rect 4893 2601 4905 2604
rect 4939 2601 4951 2635
rect 4893 2595 4951 2601
rect 6362 2592 6368 2644
rect 6420 2632 6426 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 6420 2604 6745 2632
rect 6420 2592 6426 2604
rect 6733 2601 6745 2604
rect 6779 2601 6791 2635
rect 6733 2595 6791 2601
rect 7009 2635 7067 2641
rect 7009 2601 7021 2635
rect 7055 2632 7067 2635
rect 7098 2632 7104 2644
rect 7055 2604 7104 2632
rect 7055 2601 7067 2604
rect 7009 2595 7067 2601
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7926 2592 7932 2644
rect 7984 2592 7990 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8386 2632 8392 2644
rect 8067 2604 8392 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 10502 2592 10508 2644
rect 10560 2592 10566 2644
rect 12250 2592 12256 2644
rect 12308 2632 12314 2644
rect 12345 2635 12403 2641
rect 12345 2632 12357 2635
rect 12308 2604 12357 2632
rect 12308 2592 12314 2604
rect 12345 2601 12357 2604
rect 12391 2601 12403 2635
rect 12345 2595 12403 2601
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 12492 2604 12633 2632
rect 12492 2592 12498 2604
rect 12621 2601 12633 2604
rect 12667 2601 12679 2635
rect 12621 2595 12679 2601
rect 16114 2592 16120 2644
rect 16172 2592 16178 2644
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 3896 2564 3924 2592
rect 1627 2536 3924 2564
rect 3988 2536 5488 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 2590 2456 2596 2508
rect 2648 2496 2654 2508
rect 3513 2499 3571 2505
rect 3513 2496 3525 2499
rect 2648 2468 3525 2496
rect 2648 2456 2654 2468
rect 3513 2465 3525 2468
rect 3559 2496 3571 2499
rect 3988 2496 4016 2536
rect 3559 2468 4016 2496
rect 3559 2465 3571 2468
rect 3513 2459 3571 2465
rect 4246 2456 4252 2508
rect 4304 2456 4310 2508
rect 5460 2505 5488 2536
rect 5445 2499 5503 2505
rect 5445 2465 5457 2499
rect 5491 2465 5503 2499
rect 7944 2496 7972 2592
rect 11698 2524 11704 2576
rect 11756 2564 11762 2576
rect 15841 2567 15899 2573
rect 15841 2564 15853 2567
rect 11756 2536 15853 2564
rect 11756 2524 11762 2536
rect 5445 2459 5503 2465
rect 7208 2468 7972 2496
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2428 3387 2431
rect 4264 2428 4292 2456
rect 3375 2400 4292 2428
rect 3375 2397 3387 2400
rect 3329 2391 3387 2397
rect 5350 2388 5356 2440
rect 5408 2388 5414 2440
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 7208 2437 7236 2468
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6512 2400 6561 2428
rect 6512 2388 6518 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 9953 2431 10011 2437
rect 9953 2397 9965 2431
rect 9999 2428 10011 2431
rect 10042 2428 10048 2440
rect 9999 2400 10048 2428
rect 9999 2397 10011 2400
rect 9953 2391 10011 2397
rect 3237 2363 3295 2369
rect 3237 2329 3249 2363
rect 3283 2360 3295 2363
rect 3786 2360 3792 2372
rect 3283 2332 3792 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 3786 2320 3792 2332
rect 3844 2320 3850 2372
rect 4062 2320 4068 2372
rect 4120 2320 4126 2372
rect 5261 2363 5319 2369
rect 5261 2329 5273 2363
rect 5307 2360 5319 2363
rect 5736 2360 5764 2388
rect 9968 2360 9996 2391
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 11808 2437 11836 2536
rect 15841 2533 15853 2536
rect 15887 2533 15899 2567
rect 15841 2527 15899 2533
rect 11974 2456 11980 2508
rect 12032 2496 12038 2508
rect 12032 2468 12480 2496
rect 12032 2456 12038 2468
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 11793 2431 11851 2437
rect 10367 2400 11744 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 5307 2332 5764 2360
rect 5828 2332 9996 2360
rect 10137 2363 10195 2369
rect 5307 2329 5319 2332
rect 5261 2323 5319 2329
rect 4157 2295 4215 2301
rect 4157 2261 4169 2295
rect 4203 2292 4215 2295
rect 5166 2292 5172 2304
rect 4203 2264 5172 2292
rect 4203 2261 4215 2264
rect 4157 2255 4215 2261
rect 5166 2252 5172 2264
rect 5224 2292 5230 2304
rect 5828 2292 5856 2332
rect 10137 2329 10149 2363
rect 10183 2329 10195 2363
rect 10137 2323 10195 2329
rect 10229 2363 10287 2369
rect 10229 2329 10241 2363
rect 10275 2360 10287 2363
rect 10410 2360 10416 2372
rect 10275 2332 10416 2360
rect 10275 2329 10287 2332
rect 10229 2323 10287 2329
rect 5224 2264 5856 2292
rect 10152 2292 10180 2323
rect 10410 2320 10416 2332
rect 10468 2320 10474 2372
rect 11716 2360 11744 2400
rect 11793 2397 11805 2431
rect 11839 2397 11851 2431
rect 12158 2428 12164 2440
rect 11793 2391 11851 2397
rect 11900 2400 12164 2428
rect 11900 2360 11928 2400
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 12452 2437 12480 2468
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 16347 2400 16436 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 11716 2332 11928 2360
rect 11977 2363 12035 2369
rect 11977 2329 11989 2363
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 12069 2363 12127 2369
rect 12069 2329 12081 2363
rect 12115 2360 12127 2363
rect 13354 2360 13360 2372
rect 12115 2332 13360 2360
rect 12115 2329 12127 2332
rect 12069 2323 12127 2329
rect 11790 2292 11796 2304
rect 10152 2264 11796 2292
rect 5224 2252 5230 2264
rect 11790 2252 11796 2264
rect 11848 2292 11854 2304
rect 11992 2292 12020 2323
rect 13354 2320 13360 2332
rect 13412 2320 13418 2372
rect 15654 2320 15660 2372
rect 15712 2320 15718 2372
rect 16408 2304 16436 2400
rect 11848 2264 12020 2292
rect 11848 2252 11854 2264
rect 16390 2252 16396 2304
rect 16448 2252 16454 2304
rect 1104 2202 16811 2224
rect 1104 2150 4836 2202
rect 4888 2150 4900 2202
rect 4952 2150 4964 2202
rect 5016 2150 5028 2202
rect 5080 2150 5092 2202
rect 5144 2150 8723 2202
rect 8775 2150 8787 2202
rect 8839 2150 8851 2202
rect 8903 2150 8915 2202
rect 8967 2150 8979 2202
rect 9031 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 16497 2202
rect 16549 2150 16561 2202
rect 16613 2150 16625 2202
rect 16677 2150 16689 2202
rect 16741 2150 16753 2202
rect 16805 2150 16811 2202
rect 1104 2128 16811 2150
<< via1 >>
rect 4836 17382 4888 17434
rect 4900 17382 4952 17434
rect 4964 17382 5016 17434
rect 5028 17382 5080 17434
rect 5092 17382 5144 17434
rect 8723 17382 8775 17434
rect 8787 17382 8839 17434
rect 8851 17382 8903 17434
rect 8915 17382 8967 17434
rect 8979 17382 9031 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 16497 17382 16549 17434
rect 16561 17382 16613 17434
rect 16625 17382 16677 17434
rect 16689 17382 16741 17434
rect 16753 17382 16805 17434
rect 20 17280 72 17332
rect 4620 17280 4672 17332
rect 15476 17280 15528 17332
rect 3608 17212 3660 17264
rect 7748 17212 7800 17264
rect 11612 17212 11664 17264
rect 1492 17187 1544 17196
rect 1492 17153 1501 17187
rect 1501 17153 1535 17187
rect 1535 17153 1544 17187
rect 1492 17144 1544 17153
rect 3884 17144 3936 17196
rect 7104 17144 7156 17196
rect 9312 17187 9364 17196
rect 9312 17153 9321 17187
rect 9321 17153 9355 17187
rect 9355 17153 9364 17187
rect 9312 17144 9364 17153
rect 15936 17255 15988 17264
rect 15936 17221 15945 17255
rect 15945 17221 15979 17255
rect 15979 17221 15988 17255
rect 15936 17212 15988 17221
rect 3792 17119 3844 17128
rect 3792 17085 3801 17119
rect 3801 17085 3835 17119
rect 3835 17085 3844 17119
rect 3792 17076 3844 17085
rect 9404 17119 9456 17128
rect 9404 17085 9413 17119
rect 9413 17085 9447 17119
rect 9447 17085 9456 17119
rect 9404 17076 9456 17085
rect 8300 17008 8352 17060
rect 10140 17008 10192 17060
rect 3332 16940 3384 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 8024 16983 8076 16992
rect 8024 16949 8033 16983
rect 8033 16949 8067 16983
rect 8067 16949 8076 16983
rect 8024 16940 8076 16949
rect 8116 16940 8168 16992
rect 11888 16983 11940 16992
rect 11888 16949 11897 16983
rect 11897 16949 11931 16983
rect 11931 16949 11940 16983
rect 11888 16940 11940 16949
rect 15752 16983 15804 16992
rect 15752 16949 15761 16983
rect 15761 16949 15795 16983
rect 15795 16949 15804 16983
rect 15752 16940 15804 16949
rect 2893 16838 2945 16890
rect 2957 16838 3009 16890
rect 3021 16838 3073 16890
rect 3085 16838 3137 16890
rect 3149 16838 3201 16890
rect 6780 16838 6832 16890
rect 6844 16838 6896 16890
rect 6908 16838 6960 16890
rect 6972 16838 7024 16890
rect 7036 16838 7088 16890
rect 10667 16838 10719 16890
rect 10731 16838 10783 16890
rect 10795 16838 10847 16890
rect 10859 16838 10911 16890
rect 10923 16838 10975 16890
rect 14554 16838 14606 16890
rect 14618 16838 14670 16890
rect 14682 16838 14734 16890
rect 14746 16838 14798 16890
rect 14810 16838 14862 16890
rect 3240 16736 3292 16788
rect 3884 16779 3936 16788
rect 3884 16745 3893 16779
rect 3893 16745 3927 16779
rect 3927 16745 3936 16779
rect 3884 16736 3936 16745
rect 3792 16668 3844 16720
rect 4160 16600 4212 16652
rect 6460 16600 6512 16652
rect 7104 16736 7156 16788
rect 9312 16736 9364 16788
rect 940 16532 992 16584
rect 2136 16464 2188 16516
rect 2688 16396 2740 16448
rect 2780 16396 2832 16448
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 8392 16532 8444 16584
rect 11060 16600 11112 16652
rect 6736 16464 6788 16516
rect 7288 16507 7340 16516
rect 7288 16473 7297 16507
rect 7297 16473 7331 16507
rect 7331 16473 7340 16507
rect 7288 16464 7340 16473
rect 9772 16464 9824 16516
rect 5172 16396 5224 16448
rect 9404 16396 9456 16448
rect 4836 16294 4888 16346
rect 4900 16294 4952 16346
rect 4964 16294 5016 16346
rect 5028 16294 5080 16346
rect 5092 16294 5144 16346
rect 8723 16294 8775 16346
rect 8787 16294 8839 16346
rect 8851 16294 8903 16346
rect 8915 16294 8967 16346
rect 8979 16294 9031 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 16497 16294 16549 16346
rect 16561 16294 16613 16346
rect 16625 16294 16677 16346
rect 16689 16294 16741 16346
rect 16753 16294 16805 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 2688 16192 2740 16244
rect 6276 16124 6328 16176
rect 2780 16056 2832 16108
rect 3700 16056 3752 16108
rect 3424 16031 3476 16040
rect 3424 15997 3433 16031
rect 3433 15997 3467 16031
rect 3467 15997 3476 16031
rect 3424 15988 3476 15997
rect 3792 15988 3844 16040
rect 4160 15988 4212 16040
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 6184 15852 6236 15861
rect 6460 16235 6512 16244
rect 6460 16201 6469 16235
rect 6469 16201 6503 16235
rect 6503 16201 6512 16235
rect 6460 16192 6512 16201
rect 6736 16192 6788 16244
rect 7288 16192 7340 16244
rect 8116 16192 8168 16244
rect 8392 16235 8444 16244
rect 8392 16201 8401 16235
rect 8401 16201 8435 16235
rect 8435 16201 8444 16235
rect 8392 16192 8444 16201
rect 9404 16192 9456 16244
rect 9772 16235 9824 16244
rect 9772 16201 9781 16235
rect 9781 16201 9815 16235
rect 9815 16201 9824 16235
rect 9772 16192 9824 16201
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 7932 16056 7984 16108
rect 12256 16124 12308 16176
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 10416 16056 10468 16108
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 11520 16031 11572 16040
rect 11520 15997 11529 16031
rect 11529 15997 11563 16031
rect 11563 15997 11572 16031
rect 11520 15988 11572 15997
rect 13176 15988 13228 16040
rect 13728 15920 13780 15972
rect 8392 15852 8444 15904
rect 13360 15895 13412 15904
rect 13360 15861 13369 15895
rect 13369 15861 13403 15895
rect 13403 15861 13412 15895
rect 13360 15852 13412 15861
rect 2893 15750 2945 15802
rect 2957 15750 3009 15802
rect 3021 15750 3073 15802
rect 3085 15750 3137 15802
rect 3149 15750 3201 15802
rect 6780 15750 6832 15802
rect 6844 15750 6896 15802
rect 6908 15750 6960 15802
rect 6972 15750 7024 15802
rect 7036 15750 7088 15802
rect 10667 15750 10719 15802
rect 10731 15750 10783 15802
rect 10795 15750 10847 15802
rect 10859 15750 10911 15802
rect 10923 15750 10975 15802
rect 14554 15750 14606 15802
rect 14618 15750 14670 15802
rect 14682 15750 14734 15802
rect 14746 15750 14798 15802
rect 14810 15750 14862 15802
rect 3424 15648 3476 15700
rect 4712 15648 4764 15700
rect 6276 15691 6328 15700
rect 6276 15657 6285 15691
rect 6285 15657 6319 15691
rect 6319 15657 6328 15691
rect 6276 15648 6328 15657
rect 9404 15691 9456 15700
rect 9404 15657 9413 15691
rect 9413 15657 9447 15691
rect 9447 15657 9456 15691
rect 9404 15648 9456 15657
rect 12256 15691 12308 15700
rect 12256 15657 12265 15691
rect 12265 15657 12299 15691
rect 12299 15657 12308 15691
rect 12256 15648 12308 15657
rect 13360 15648 13412 15700
rect 5172 15623 5224 15632
rect 5172 15589 5181 15623
rect 5181 15589 5215 15623
rect 5215 15589 5224 15623
rect 5172 15580 5224 15589
rect 10232 15580 10284 15632
rect 11888 15580 11940 15632
rect 3700 15444 3752 15496
rect 4896 15487 4948 15496
rect 4896 15453 4905 15487
rect 4905 15453 4939 15487
rect 4939 15453 4948 15487
rect 4896 15444 4948 15453
rect 5264 15444 5316 15496
rect 7932 15444 7984 15496
rect 4896 15308 4948 15360
rect 5448 15308 5500 15360
rect 8024 15308 8076 15360
rect 9220 15308 9272 15360
rect 10416 15376 10468 15428
rect 14372 15444 14424 15496
rect 10048 15308 10100 15360
rect 13084 15308 13136 15360
rect 14188 15351 14240 15360
rect 14188 15317 14197 15351
rect 14197 15317 14231 15351
rect 14231 15317 14240 15351
rect 14188 15308 14240 15317
rect 4836 15206 4888 15258
rect 4900 15206 4952 15258
rect 4964 15206 5016 15258
rect 5028 15206 5080 15258
rect 5092 15206 5144 15258
rect 8723 15206 8775 15258
rect 8787 15206 8839 15258
rect 8851 15206 8903 15258
rect 8915 15206 8967 15258
rect 8979 15206 9031 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 16497 15206 16549 15258
rect 16561 15206 16613 15258
rect 16625 15206 16677 15258
rect 16689 15206 16741 15258
rect 16753 15206 16805 15258
rect 1492 15104 1544 15156
rect 2320 15104 2372 15156
rect 7656 15104 7708 15156
rect 8300 15104 8352 15156
rect 1676 15011 1728 15020
rect 1676 14977 1710 15011
rect 1710 14977 1728 15011
rect 1676 14968 1728 14977
rect 7748 15011 7800 15020
rect 7748 14977 7757 15011
rect 7757 14977 7791 15011
rect 7791 14977 7800 15011
rect 7748 14968 7800 14977
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 9128 15036 9180 15088
rect 9312 15036 9364 15088
rect 10508 15036 10560 15088
rect 11520 15036 11572 15088
rect 12256 15036 12308 15088
rect 8576 14832 8628 14884
rect 7472 14764 7524 14816
rect 13084 15036 13136 15088
rect 14188 15036 14240 15088
rect 9864 14943 9916 14952
rect 9864 14909 9873 14943
rect 9873 14909 9907 14943
rect 9907 14909 9916 14943
rect 9864 14900 9916 14909
rect 11244 14900 11296 14952
rect 11336 14900 11388 14952
rect 11980 14943 12032 14952
rect 11980 14909 11989 14943
rect 11989 14909 12023 14943
rect 12023 14909 12032 14943
rect 11980 14900 12032 14909
rect 13728 14900 13780 14952
rect 13636 14764 13688 14816
rect 14464 14764 14516 14816
rect 2893 14662 2945 14714
rect 2957 14662 3009 14714
rect 3021 14662 3073 14714
rect 3085 14662 3137 14714
rect 3149 14662 3201 14714
rect 6780 14662 6832 14714
rect 6844 14662 6896 14714
rect 6908 14662 6960 14714
rect 6972 14662 7024 14714
rect 7036 14662 7088 14714
rect 10667 14662 10719 14714
rect 10731 14662 10783 14714
rect 10795 14662 10847 14714
rect 10859 14662 10911 14714
rect 10923 14662 10975 14714
rect 14554 14662 14606 14714
rect 14618 14662 14670 14714
rect 14682 14662 14734 14714
rect 14746 14662 14798 14714
rect 14810 14662 14862 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 1400 14424 1452 14476
rect 5172 14535 5224 14544
rect 5172 14501 5181 14535
rect 5181 14501 5215 14535
rect 5215 14501 5224 14535
rect 5172 14492 5224 14501
rect 7748 14560 7800 14612
rect 9864 14560 9916 14612
rect 10508 14560 10560 14612
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 3792 14467 3844 14476
rect 3792 14433 3801 14467
rect 3801 14433 3835 14467
rect 3835 14433 3844 14467
rect 3792 14424 3844 14433
rect 8300 14492 8352 14544
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 3332 14399 3384 14408
rect 3332 14365 3341 14399
rect 3341 14365 3375 14399
rect 3375 14365 3384 14399
rect 3332 14356 3384 14365
rect 3700 14356 3752 14408
rect 4896 14356 4948 14408
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 7656 14356 7708 14408
rect 7932 14356 7984 14408
rect 10416 14492 10468 14544
rect 9588 14467 9640 14476
rect 9588 14433 9597 14467
rect 9597 14433 9631 14467
rect 9631 14433 9640 14467
rect 9588 14424 9640 14433
rect 9404 14399 9456 14408
rect 9404 14365 9413 14399
rect 9413 14365 9447 14399
rect 9447 14365 9456 14399
rect 9404 14356 9456 14365
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 11060 14424 11112 14476
rect 13728 14424 13780 14476
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 14464 14356 14516 14365
rect 2596 14220 2648 14272
rect 3608 14263 3660 14272
rect 3608 14229 3617 14263
rect 3617 14229 3651 14263
rect 3651 14229 3660 14263
rect 3608 14220 3660 14229
rect 3884 14220 3936 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 8576 14288 8628 14340
rect 11520 14288 11572 14340
rect 12348 14288 12400 14340
rect 10508 14220 10560 14272
rect 14096 14263 14148 14272
rect 14096 14229 14105 14263
rect 14105 14229 14139 14263
rect 14139 14229 14148 14263
rect 14096 14220 14148 14229
rect 14280 14220 14332 14272
rect 16212 14220 16264 14272
rect 4836 14118 4888 14170
rect 4900 14118 4952 14170
rect 4964 14118 5016 14170
rect 5028 14118 5080 14170
rect 5092 14118 5144 14170
rect 8723 14118 8775 14170
rect 8787 14118 8839 14170
rect 8851 14118 8903 14170
rect 8915 14118 8967 14170
rect 8979 14118 9031 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 16497 14118 16549 14170
rect 16561 14118 16613 14170
rect 16625 14118 16677 14170
rect 16689 14118 16741 14170
rect 16753 14118 16805 14170
rect 1768 14016 1820 14068
rect 2780 14016 2832 14068
rect 3148 14016 3200 14068
rect 3608 14016 3660 14068
rect 4712 14016 4764 14068
rect 5172 14016 5224 14068
rect 7840 14016 7892 14068
rect 8576 14016 8628 14068
rect 9404 14016 9456 14068
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 12348 14059 12400 14068
rect 12348 14025 12357 14059
rect 12357 14025 12391 14059
rect 12391 14025 12400 14059
rect 12348 14016 12400 14025
rect 13176 14016 13228 14068
rect 14096 14016 14148 14068
rect 14372 14016 14424 14068
rect 16212 14059 16264 14068
rect 16212 14025 16221 14059
rect 16221 14025 16255 14059
rect 16255 14025 16264 14059
rect 16212 14016 16264 14025
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 3424 13812 3476 13864
rect 3884 13812 3936 13864
rect 4068 13855 4120 13864
rect 4068 13821 4077 13855
rect 4077 13821 4111 13855
rect 4111 13821 4120 13855
rect 4068 13812 4120 13821
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 5632 13880 5684 13932
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 11428 13948 11480 14000
rect 10324 13923 10376 13932
rect 10324 13889 10333 13923
rect 10333 13889 10367 13923
rect 10367 13889 10376 13923
rect 10324 13880 10376 13889
rect 11060 13880 11112 13932
rect 11520 13880 11572 13932
rect 5264 13855 5316 13864
rect 5264 13821 5273 13855
rect 5273 13821 5307 13855
rect 5307 13821 5316 13855
rect 5264 13812 5316 13821
rect 9220 13812 9272 13864
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 12992 13880 13044 13932
rect 9128 13744 9180 13796
rect 12072 13812 12124 13864
rect 12256 13812 12308 13864
rect 15384 13948 15436 14000
rect 11244 13744 11296 13796
rect 5632 13676 5684 13728
rect 16580 13812 16632 13864
rect 14372 13744 14424 13796
rect 13820 13676 13872 13728
rect 14280 13719 14332 13728
rect 14280 13685 14289 13719
rect 14289 13685 14323 13719
rect 14323 13685 14332 13719
rect 14280 13676 14332 13685
rect 2893 13574 2945 13626
rect 2957 13574 3009 13626
rect 3021 13574 3073 13626
rect 3085 13574 3137 13626
rect 3149 13574 3201 13626
rect 6780 13574 6832 13626
rect 6844 13574 6896 13626
rect 6908 13574 6960 13626
rect 6972 13574 7024 13626
rect 7036 13574 7088 13626
rect 10667 13574 10719 13626
rect 10731 13574 10783 13626
rect 10795 13574 10847 13626
rect 10859 13574 10911 13626
rect 10923 13574 10975 13626
rect 14554 13574 14606 13626
rect 14618 13574 14670 13626
rect 14682 13574 14734 13626
rect 14746 13574 14798 13626
rect 14810 13574 14862 13626
rect 5264 13472 5316 13524
rect 10324 13472 10376 13524
rect 11060 13472 11112 13524
rect 12992 13472 13044 13524
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 5632 13336 5684 13388
rect 9312 13336 9364 13388
rect 13820 13336 13872 13388
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 6184 13268 6236 13320
rect 7288 13268 7340 13320
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 3056 13175 3108 13184
rect 3056 13141 3065 13175
rect 3065 13141 3099 13175
rect 3099 13141 3108 13175
rect 3056 13132 3108 13141
rect 3332 13132 3384 13184
rect 9496 13200 9548 13252
rect 9956 13132 10008 13184
rect 11428 13268 11480 13320
rect 11336 13200 11388 13252
rect 11888 13200 11940 13252
rect 12164 13200 12216 13252
rect 11152 13132 11204 13184
rect 12440 13132 12492 13184
rect 14280 13200 14332 13252
rect 15384 13200 15436 13252
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 4836 13030 4888 13082
rect 4900 13030 4952 13082
rect 4964 13030 5016 13082
rect 5028 13030 5080 13082
rect 5092 13030 5144 13082
rect 8723 13030 8775 13082
rect 8787 13030 8839 13082
rect 8851 13030 8903 13082
rect 8915 13030 8967 13082
rect 8979 13030 9031 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 16497 13030 16549 13082
rect 16561 13030 16613 13082
rect 16625 13030 16677 13082
rect 16689 13030 16741 13082
rect 16753 13030 16805 13082
rect 4712 12928 4764 12980
rect 6184 12928 6236 12980
rect 8300 12928 8352 12980
rect 4160 12860 4212 12912
rect 7104 12860 7156 12912
rect 8576 12903 8628 12912
rect 8576 12869 8585 12903
rect 8585 12869 8619 12903
rect 8619 12869 8628 12903
rect 8576 12860 8628 12869
rect 2320 12835 2372 12844
rect 2320 12801 2329 12835
rect 2329 12801 2363 12835
rect 2363 12801 2372 12835
rect 2320 12792 2372 12801
rect 2688 12792 2740 12844
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 3516 12724 3568 12776
rect 5908 12767 5960 12776
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2780 12588 2832 12640
rect 5724 12588 5776 12640
rect 6368 12767 6420 12776
rect 6368 12733 6377 12767
rect 6377 12733 6411 12767
rect 6411 12733 6420 12767
rect 6368 12724 6420 12733
rect 6644 12767 6696 12776
rect 6644 12733 6653 12767
rect 6653 12733 6687 12767
rect 6687 12733 6696 12767
rect 6644 12724 6696 12733
rect 7932 12724 7984 12776
rect 9128 12928 9180 12980
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 10232 12928 10284 12980
rect 10416 12860 10468 12912
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 11060 12903 11112 12912
rect 11060 12869 11069 12903
rect 11069 12869 11103 12903
rect 11103 12869 11112 12903
rect 11060 12860 11112 12869
rect 11336 12971 11388 12980
rect 11336 12937 11345 12971
rect 11345 12937 11379 12971
rect 11379 12937 11388 12971
rect 11336 12928 11388 12937
rect 11796 12860 11848 12912
rect 12072 12860 12124 12912
rect 12440 12928 12492 12980
rect 15844 12928 15896 12980
rect 13360 12903 13412 12912
rect 13360 12869 13369 12903
rect 13369 12869 13403 12903
rect 13403 12869 13412 12903
rect 13360 12860 13412 12869
rect 11888 12792 11940 12844
rect 8668 12656 8720 12708
rect 8116 12631 8168 12640
rect 8116 12597 8125 12631
rect 8125 12597 8159 12631
rect 8159 12597 8168 12631
rect 8116 12588 8168 12597
rect 8392 12588 8444 12640
rect 10048 12588 10100 12640
rect 12164 12724 12216 12776
rect 13728 12860 13780 12912
rect 13820 12860 13872 12912
rect 13636 12792 13688 12844
rect 13912 12724 13964 12776
rect 12532 12631 12584 12640
rect 12532 12597 12541 12631
rect 12541 12597 12575 12631
rect 12575 12597 12584 12631
rect 12532 12588 12584 12597
rect 13820 12588 13872 12640
rect 2893 12486 2945 12538
rect 2957 12486 3009 12538
rect 3021 12486 3073 12538
rect 3085 12486 3137 12538
rect 3149 12486 3201 12538
rect 6780 12486 6832 12538
rect 6844 12486 6896 12538
rect 6908 12486 6960 12538
rect 6972 12486 7024 12538
rect 7036 12486 7088 12538
rect 10667 12486 10719 12538
rect 10731 12486 10783 12538
rect 10795 12486 10847 12538
rect 10859 12486 10911 12538
rect 10923 12486 10975 12538
rect 14554 12486 14606 12538
rect 14618 12486 14670 12538
rect 14682 12486 14734 12538
rect 14746 12486 14798 12538
rect 14810 12486 14862 12538
rect 2044 12384 2096 12436
rect 3240 12384 3292 12436
rect 4160 12384 4212 12436
rect 5356 12384 5408 12436
rect 6644 12384 6696 12436
rect 7104 12384 7156 12436
rect 7288 12427 7340 12436
rect 7288 12393 7297 12427
rect 7297 12393 7331 12427
rect 7331 12393 7340 12427
rect 7288 12384 7340 12393
rect 8484 12384 8536 12436
rect 2688 12316 2740 12368
rect 1768 12248 1820 12300
rect 2320 12248 2372 12300
rect 5540 12248 5592 12300
rect 7932 12291 7984 12300
rect 7932 12257 7941 12291
rect 7941 12257 7975 12291
rect 7975 12257 7984 12291
rect 7932 12248 7984 12257
rect 11980 12384 12032 12436
rect 13360 12384 13412 12436
rect 2780 12180 2832 12232
rect 3884 12223 3936 12232
rect 3884 12189 3893 12223
rect 3893 12189 3927 12223
rect 3927 12189 3936 12223
rect 3884 12180 3936 12189
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 7656 12180 7708 12232
rect 9772 12180 9824 12232
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 8116 12112 8168 12164
rect 9312 12112 9364 12164
rect 12072 12112 12124 12164
rect 12532 12223 12584 12232
rect 12532 12189 12566 12223
rect 12566 12189 12584 12223
rect 12532 12180 12584 12189
rect 13820 12180 13872 12232
rect 15752 12112 15804 12164
rect 7932 12044 7984 12096
rect 10232 12044 10284 12096
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 4836 11942 4888 11994
rect 4900 11942 4952 11994
rect 4964 11942 5016 11994
rect 5028 11942 5080 11994
rect 5092 11942 5144 11994
rect 8723 11942 8775 11994
rect 8787 11942 8839 11994
rect 8851 11942 8903 11994
rect 8915 11942 8967 11994
rect 8979 11942 9031 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 16497 11942 16549 11994
rect 16561 11942 16613 11994
rect 16625 11942 16677 11994
rect 16689 11942 16741 11994
rect 16753 11942 16805 11994
rect 3976 11840 4028 11892
rect 9312 11840 9364 11892
rect 12072 11883 12124 11892
rect 12072 11849 12081 11883
rect 12081 11849 12115 11883
rect 12115 11849 12124 11883
rect 12072 11840 12124 11849
rect 14096 11840 14148 11892
rect 2780 11704 2832 11756
rect 6368 11704 6420 11756
rect 6644 11704 6696 11756
rect 8024 11772 8076 11824
rect 11704 11815 11756 11824
rect 11704 11781 11713 11815
rect 11713 11781 11747 11815
rect 11747 11781 11756 11815
rect 11704 11772 11756 11781
rect 11980 11772 12032 11824
rect 15016 11772 15068 11824
rect 9404 11747 9456 11756
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 11336 11704 11388 11756
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 12256 11704 12308 11756
rect 15844 11636 15896 11688
rect 1860 11500 1912 11552
rect 2228 11500 2280 11552
rect 3884 11500 3936 11552
rect 9772 11568 9824 11620
rect 10232 11568 10284 11620
rect 7932 11543 7984 11552
rect 7932 11509 7941 11543
rect 7941 11509 7975 11543
rect 7975 11509 7984 11543
rect 7932 11500 7984 11509
rect 8300 11500 8352 11552
rect 9588 11500 9640 11552
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 2893 11398 2945 11450
rect 2957 11398 3009 11450
rect 3021 11398 3073 11450
rect 3085 11398 3137 11450
rect 3149 11398 3201 11450
rect 6780 11398 6832 11450
rect 6844 11398 6896 11450
rect 6908 11398 6960 11450
rect 6972 11398 7024 11450
rect 7036 11398 7088 11450
rect 10667 11398 10719 11450
rect 10731 11398 10783 11450
rect 10795 11398 10847 11450
rect 10859 11398 10911 11450
rect 10923 11398 10975 11450
rect 14554 11398 14606 11450
rect 14618 11398 14670 11450
rect 14682 11398 14734 11450
rect 14746 11398 14798 11450
rect 14810 11398 14862 11450
rect 3332 11339 3384 11348
rect 3332 11305 3341 11339
rect 3341 11305 3375 11339
rect 3375 11305 3384 11339
rect 3332 11296 3384 11305
rect 4068 11296 4120 11348
rect 3976 11228 4028 11280
rect 3792 11203 3844 11212
rect 3792 11169 3801 11203
rect 3801 11169 3835 11203
rect 3835 11169 3844 11203
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 8208 11296 8260 11348
rect 8668 11296 8720 11348
rect 9036 11296 9088 11348
rect 9404 11296 9456 11348
rect 6092 11271 6144 11280
rect 6092 11237 6101 11271
rect 6101 11237 6135 11271
rect 6135 11237 6144 11271
rect 6092 11228 6144 11237
rect 3792 11160 3844 11169
rect 8300 11228 8352 11280
rect 9220 11228 9272 11280
rect 1860 11135 1912 11144
rect 1860 11101 1869 11135
rect 1869 11101 1903 11135
rect 1903 11101 1912 11135
rect 1860 11092 1912 11101
rect 2044 11092 2096 11144
rect 2228 11135 2280 11144
rect 2228 11101 2262 11135
rect 2262 11101 2280 11135
rect 2228 11092 2280 11101
rect 3700 11092 3752 11144
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 4160 10999 4212 11008
rect 4160 10965 4169 10999
rect 4169 10965 4203 10999
rect 4203 10965 4212 10999
rect 4160 10956 4212 10965
rect 6000 11092 6052 11144
rect 7932 11092 7984 11144
rect 4712 11024 4764 11076
rect 5816 11024 5868 11076
rect 8484 11160 8536 11212
rect 8576 11160 8628 11212
rect 14280 11296 14332 11348
rect 15476 11296 15528 11348
rect 15844 11339 15896 11348
rect 15844 11305 15853 11339
rect 15853 11305 15887 11339
rect 15887 11305 15896 11339
rect 15844 11296 15896 11305
rect 9772 11092 9824 11144
rect 9864 11092 9916 11144
rect 10508 11092 10560 11144
rect 11888 11160 11940 11212
rect 15200 11228 15252 11280
rect 9404 11024 9456 11076
rect 9956 11024 10008 11076
rect 11704 11092 11756 11144
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 14924 11203 14976 11212
rect 14924 11169 14933 11203
rect 14933 11169 14967 11203
rect 14967 11169 14976 11203
rect 14924 11160 14976 11169
rect 15752 11271 15804 11280
rect 15752 11237 15761 11271
rect 15761 11237 15795 11271
rect 15795 11237 15804 11271
rect 15752 11228 15804 11237
rect 16120 11024 16172 11076
rect 6368 10956 6420 11008
rect 7012 10999 7064 11008
rect 7012 10965 7021 10999
rect 7021 10965 7055 10999
rect 7055 10965 7064 10999
rect 7012 10956 7064 10965
rect 7472 10999 7524 11008
rect 7472 10965 7481 10999
rect 7481 10965 7515 10999
rect 7515 10965 7524 10999
rect 7472 10956 7524 10965
rect 8484 10956 8536 11008
rect 4836 10854 4888 10906
rect 4900 10854 4952 10906
rect 4964 10854 5016 10906
rect 5028 10854 5080 10906
rect 5092 10854 5144 10906
rect 8723 10854 8775 10906
rect 8787 10854 8839 10906
rect 8851 10854 8903 10906
rect 8915 10854 8967 10906
rect 8979 10854 9031 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 16497 10854 16549 10906
rect 16561 10854 16613 10906
rect 16625 10854 16677 10906
rect 16689 10854 16741 10906
rect 16753 10854 16805 10906
rect 2780 10752 2832 10804
rect 3332 10752 3384 10804
rect 4160 10752 4212 10804
rect 4712 10752 4764 10804
rect 5816 10795 5868 10804
rect 5816 10761 5825 10795
rect 5825 10761 5859 10795
rect 5859 10761 5868 10795
rect 5816 10752 5868 10761
rect 6092 10752 6144 10804
rect 6644 10752 6696 10804
rect 7012 10752 7064 10804
rect 7472 10795 7524 10804
rect 7472 10761 7481 10795
rect 7481 10761 7515 10795
rect 7515 10761 7524 10795
rect 7472 10752 7524 10761
rect 8484 10752 8536 10804
rect 9404 10752 9456 10804
rect 9496 10752 9548 10804
rect 9772 10752 9824 10804
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 12072 10752 12124 10804
rect 14280 10752 14332 10804
rect 15016 10752 15068 10804
rect 15200 10752 15252 10804
rect 1676 10727 1728 10736
rect 1676 10693 1710 10727
rect 1710 10693 1728 10727
rect 1676 10684 1728 10693
rect 2044 10616 2096 10668
rect 3700 10616 3752 10668
rect 3884 10616 3936 10668
rect 8300 10684 8352 10736
rect 3516 10412 3568 10464
rect 4344 10591 4396 10600
rect 4344 10557 4353 10591
rect 4353 10557 4387 10591
rect 4387 10557 4396 10591
rect 4344 10548 4396 10557
rect 5356 10548 5408 10600
rect 7196 10548 7248 10600
rect 8116 10548 8168 10600
rect 8576 10548 8628 10600
rect 8300 10480 8352 10532
rect 9128 10548 9180 10600
rect 9680 10684 9732 10736
rect 10600 10684 10652 10736
rect 9496 10548 9548 10600
rect 10140 10616 10192 10668
rect 11060 10659 11112 10668
rect 9772 10591 9824 10600
rect 9772 10557 9781 10591
rect 9781 10557 9815 10591
rect 9815 10557 9824 10591
rect 9772 10548 9824 10557
rect 11060 10625 11069 10659
rect 11069 10625 11103 10659
rect 11103 10625 11112 10659
rect 11060 10616 11112 10625
rect 13912 10616 13964 10668
rect 14280 10616 14332 10668
rect 15016 10616 15068 10668
rect 4068 10412 4120 10464
rect 8392 10412 8444 10464
rect 9772 10412 9824 10464
rect 10140 10412 10192 10464
rect 13728 10412 13780 10464
rect 15108 10455 15160 10464
rect 15108 10421 15117 10455
rect 15117 10421 15151 10455
rect 15151 10421 15160 10455
rect 15108 10412 15160 10421
rect 2893 10310 2945 10362
rect 2957 10310 3009 10362
rect 3021 10310 3073 10362
rect 3085 10310 3137 10362
rect 3149 10310 3201 10362
rect 6780 10310 6832 10362
rect 6844 10310 6896 10362
rect 6908 10310 6960 10362
rect 6972 10310 7024 10362
rect 7036 10310 7088 10362
rect 10667 10310 10719 10362
rect 10731 10310 10783 10362
rect 10795 10310 10847 10362
rect 10859 10310 10911 10362
rect 10923 10310 10975 10362
rect 14554 10310 14606 10362
rect 14618 10310 14670 10362
rect 14682 10310 14734 10362
rect 14746 10310 14798 10362
rect 14810 10310 14862 10362
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 5356 10140 5408 10192
rect 8300 10208 8352 10260
rect 9404 10208 9456 10260
rect 9680 10251 9732 10260
rect 9680 10217 9689 10251
rect 9689 10217 9723 10251
rect 9723 10217 9732 10251
rect 9680 10208 9732 10217
rect 9956 10251 10008 10260
rect 9956 10217 9965 10251
rect 9965 10217 9999 10251
rect 9999 10217 10008 10251
rect 9956 10208 10008 10217
rect 11152 10208 11204 10260
rect 11888 10208 11940 10260
rect 13912 10251 13964 10260
rect 9128 10140 9180 10192
rect 2044 10072 2096 10124
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 9956 10072 10008 10124
rect 10324 10072 10376 10124
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 5632 10004 5684 10056
rect 4528 9936 4580 9988
rect 6184 9868 6236 9920
rect 6920 9936 6972 9988
rect 9312 9936 9364 9988
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 9772 9936 9824 9988
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 9588 9868 9640 9920
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 12440 10072 12492 10124
rect 15108 10072 15160 10124
rect 13728 10004 13780 10056
rect 15384 9936 15436 9988
rect 14556 9868 14608 9920
rect 4836 9766 4888 9818
rect 4900 9766 4952 9818
rect 4964 9766 5016 9818
rect 5028 9766 5080 9818
rect 5092 9766 5144 9818
rect 8723 9766 8775 9818
rect 8787 9766 8839 9818
rect 8851 9766 8903 9818
rect 8915 9766 8967 9818
rect 8979 9766 9031 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 16497 9766 16549 9818
rect 16561 9766 16613 9818
rect 16625 9766 16677 9818
rect 16689 9766 16741 9818
rect 16753 9766 16805 9818
rect 3608 9664 3660 9716
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 6368 9664 6420 9716
rect 6920 9707 6972 9716
rect 6920 9673 6929 9707
rect 6929 9673 6963 9707
rect 6963 9673 6972 9707
rect 6920 9664 6972 9673
rect 9680 9664 9732 9716
rect 4344 9596 4396 9648
rect 1492 9528 1544 9580
rect 1676 9571 1728 9580
rect 1676 9537 1710 9571
rect 1710 9537 1728 9571
rect 1676 9528 1728 9537
rect 3884 9571 3936 9580
rect 3884 9537 3893 9571
rect 3893 9537 3927 9571
rect 3927 9537 3936 9571
rect 3884 9528 3936 9537
rect 6184 9596 6236 9648
rect 2780 9435 2832 9444
rect 2780 9401 2789 9435
rect 2789 9401 2823 9435
rect 2823 9401 2832 9435
rect 4160 9460 4212 9512
rect 6552 9528 6604 9580
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 8484 9571 8536 9580
rect 8484 9537 8493 9571
rect 8493 9537 8527 9571
rect 8527 9537 8536 9571
rect 8484 9528 8536 9537
rect 8852 9528 8904 9580
rect 12072 9664 12124 9716
rect 13912 9664 13964 9716
rect 14556 9707 14608 9716
rect 14556 9673 14565 9707
rect 14565 9673 14599 9707
rect 14599 9673 14608 9707
rect 14556 9664 14608 9673
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 8576 9460 8628 9512
rect 9496 9460 9548 9512
rect 10416 9528 10468 9580
rect 11152 9571 11204 9580
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 2780 9392 2832 9401
rect 9588 9392 9640 9444
rect 10324 9460 10376 9512
rect 15016 9596 15068 9648
rect 9312 9367 9364 9376
rect 9312 9333 9321 9367
rect 9321 9333 9355 9367
rect 9355 9333 9364 9367
rect 9312 9324 9364 9333
rect 9496 9367 9548 9376
rect 9496 9333 9505 9367
rect 9505 9333 9539 9367
rect 9539 9333 9548 9367
rect 9496 9324 9548 9333
rect 10232 9367 10284 9376
rect 10232 9333 10241 9367
rect 10241 9333 10275 9367
rect 10275 9333 10284 9367
rect 10232 9324 10284 9333
rect 12900 9435 12952 9444
rect 12900 9401 12909 9435
rect 12909 9401 12943 9435
rect 12943 9401 12952 9435
rect 12900 9392 12952 9401
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 14924 9460 14976 9512
rect 11888 9324 11940 9376
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 2893 9222 2945 9274
rect 2957 9222 3009 9274
rect 3021 9222 3073 9274
rect 3085 9222 3137 9274
rect 3149 9222 3201 9274
rect 6780 9222 6832 9274
rect 6844 9222 6896 9274
rect 6908 9222 6960 9274
rect 6972 9222 7024 9274
rect 7036 9222 7088 9274
rect 10667 9222 10719 9274
rect 10731 9222 10783 9274
rect 10795 9222 10847 9274
rect 10859 9222 10911 9274
rect 10923 9222 10975 9274
rect 14554 9222 14606 9274
rect 14618 9222 14670 9274
rect 14682 9222 14734 9274
rect 14746 9222 14798 9274
rect 14810 9222 14862 9274
rect 1676 9120 1728 9172
rect 2780 9120 2832 9172
rect 8484 9120 8536 9172
rect 9312 9120 9364 9172
rect 9496 9120 9548 9172
rect 9864 9120 9916 9172
rect 2596 8984 2648 9036
rect 8300 9052 8352 9104
rect 4344 8984 4396 9036
rect 5448 9027 5500 9036
rect 5448 8993 5457 9027
rect 5457 8993 5491 9027
rect 5491 8993 5500 9027
rect 5448 8984 5500 8993
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 8024 8984 8076 9036
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8484 8984 8536 9036
rect 9680 9052 9732 9104
rect 11244 9120 11296 9172
rect 12900 9120 12952 9172
rect 8852 8916 8904 8968
rect 9220 8916 9272 8968
rect 10140 8984 10192 9036
rect 11060 8984 11112 9036
rect 14924 9120 14976 9172
rect 15016 8984 15068 9036
rect 15108 8984 15160 9036
rect 10232 8916 10284 8968
rect 11520 8891 11572 8900
rect 2320 8823 2372 8832
rect 2320 8789 2329 8823
rect 2329 8789 2363 8823
rect 2363 8789 2372 8823
rect 2320 8780 2372 8789
rect 3976 8823 4028 8832
rect 3976 8789 3985 8823
rect 3985 8789 4019 8823
rect 4019 8789 4028 8823
rect 3976 8780 4028 8789
rect 5172 8823 5224 8832
rect 5172 8789 5181 8823
rect 5181 8789 5215 8823
rect 5215 8789 5224 8823
rect 5172 8780 5224 8789
rect 5816 8823 5868 8832
rect 5816 8789 5825 8823
rect 5825 8789 5859 8823
rect 5859 8789 5868 8823
rect 5816 8780 5868 8789
rect 8116 8780 8168 8832
rect 11520 8857 11529 8891
rect 11529 8857 11563 8891
rect 11563 8857 11572 8891
rect 11520 8848 11572 8857
rect 13912 8916 13964 8968
rect 8576 8780 8628 8832
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 12532 8780 12584 8832
rect 4836 8678 4888 8730
rect 4900 8678 4952 8730
rect 4964 8678 5016 8730
rect 5028 8678 5080 8730
rect 5092 8678 5144 8730
rect 8723 8678 8775 8730
rect 8787 8678 8839 8730
rect 8851 8678 8903 8730
rect 8915 8678 8967 8730
rect 8979 8678 9031 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 16497 8678 16549 8730
rect 16561 8678 16613 8730
rect 16625 8678 16677 8730
rect 16689 8678 16741 8730
rect 16753 8678 16805 8730
rect 2320 8576 2372 8628
rect 3884 8576 3936 8628
rect 5172 8576 5224 8628
rect 8484 8576 8536 8628
rect 8576 8576 8628 8628
rect 11520 8576 11572 8628
rect 12532 8576 12584 8628
rect 1492 8508 1544 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 2504 8440 2556 8492
rect 2780 8508 2832 8560
rect 3976 8440 4028 8492
rect 7196 8508 7248 8560
rect 7104 8440 7156 8492
rect 4528 8372 4580 8424
rect 9220 8440 9272 8492
rect 8208 8372 8260 8424
rect 9036 8372 9088 8424
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 9680 8440 9732 8492
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 10324 8372 10376 8424
rect 12440 8372 12492 8424
rect 9680 8304 9732 8356
rect 10416 8304 10468 8356
rect 11060 8347 11112 8356
rect 11060 8313 11069 8347
rect 11069 8313 11103 8347
rect 11103 8313 11112 8347
rect 11060 8304 11112 8313
rect 11796 8304 11848 8356
rect 6184 8279 6236 8288
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6184 8236 6236 8245
rect 6644 8236 6696 8288
rect 8484 8236 8536 8288
rect 12532 8236 12584 8288
rect 2893 8134 2945 8186
rect 2957 8134 3009 8186
rect 3021 8134 3073 8186
rect 3085 8134 3137 8186
rect 3149 8134 3201 8186
rect 6780 8134 6832 8186
rect 6844 8134 6896 8186
rect 6908 8134 6960 8186
rect 6972 8134 7024 8186
rect 7036 8134 7088 8186
rect 10667 8134 10719 8186
rect 10731 8134 10783 8186
rect 10795 8134 10847 8186
rect 10859 8134 10911 8186
rect 10923 8134 10975 8186
rect 14554 8134 14606 8186
rect 14618 8134 14670 8186
rect 14682 8134 14734 8186
rect 14746 8134 14798 8186
rect 14810 8134 14862 8186
rect 2780 8032 2832 8084
rect 5356 8075 5408 8084
rect 5356 8041 5365 8075
rect 5365 8041 5399 8075
rect 5399 8041 5408 8075
rect 5356 8032 5408 8041
rect 2596 7896 2648 7948
rect 4160 7896 4212 7948
rect 5356 7896 5408 7948
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 9404 8032 9456 8084
rect 9956 8032 10008 8084
rect 10968 8032 11020 8084
rect 11888 8032 11940 8084
rect 8484 7964 8536 8016
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 6184 7828 6236 7880
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 4068 7760 4120 7812
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 9036 7828 9088 7880
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 11060 7964 11112 8016
rect 12532 7896 12584 7948
rect 14924 7896 14976 7948
rect 10968 7828 11020 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 11980 7828 12032 7880
rect 13820 7828 13872 7880
rect 9312 7803 9364 7812
rect 9312 7769 9330 7803
rect 9330 7769 9364 7803
rect 9312 7760 9364 7769
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 6644 7692 6696 7744
rect 7380 7692 7432 7744
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 8576 7692 8628 7744
rect 9956 7803 10008 7812
rect 9956 7769 9965 7803
rect 9965 7769 9999 7803
rect 9999 7769 10008 7803
rect 9956 7760 10008 7769
rect 10232 7735 10284 7744
rect 10232 7701 10241 7735
rect 10241 7701 10275 7735
rect 10275 7701 10284 7735
rect 10232 7692 10284 7701
rect 11152 7692 11204 7744
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 13728 7760 13780 7812
rect 14096 7735 14148 7744
rect 14096 7701 14105 7735
rect 14105 7701 14139 7735
rect 14139 7701 14148 7735
rect 14096 7692 14148 7701
rect 4836 7590 4888 7642
rect 4900 7590 4952 7642
rect 4964 7590 5016 7642
rect 5028 7590 5080 7642
rect 5092 7590 5144 7642
rect 8723 7590 8775 7642
rect 8787 7590 8839 7642
rect 8851 7590 8903 7642
rect 8915 7590 8967 7642
rect 8979 7590 9031 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 16497 7590 16549 7642
rect 16561 7590 16613 7642
rect 16625 7590 16677 7642
rect 16689 7590 16741 7642
rect 16753 7590 16805 7642
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 4068 7488 4120 7540
rect 4160 7488 4212 7540
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 7104 7488 7156 7540
rect 7380 7531 7432 7540
rect 7380 7497 7389 7531
rect 7389 7497 7423 7531
rect 7423 7497 7432 7531
rect 7380 7488 7432 7497
rect 8300 7488 8352 7540
rect 10232 7488 10284 7540
rect 12072 7488 12124 7540
rect 1492 7352 1544 7404
rect 1676 7395 1728 7404
rect 1676 7361 1710 7395
rect 1710 7361 1728 7395
rect 1676 7352 1728 7361
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 13820 7488 13872 7540
rect 14096 7488 14148 7540
rect 4436 7352 4488 7404
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 5724 7352 5776 7404
rect 5908 7327 5960 7336
rect 5908 7293 5917 7327
rect 5917 7293 5951 7327
rect 5951 7293 5960 7327
rect 5908 7284 5960 7293
rect 4528 7216 4580 7268
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 8484 7148 8536 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 11060 7352 11112 7404
rect 12072 7352 12124 7404
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 15108 7420 15160 7472
rect 13636 7352 13688 7361
rect 15752 7352 15804 7404
rect 11428 7148 11480 7200
rect 11980 7148 12032 7200
rect 14004 7191 14056 7200
rect 14004 7157 14013 7191
rect 14013 7157 14047 7191
rect 14047 7157 14056 7191
rect 14004 7148 14056 7157
rect 15384 7148 15436 7200
rect 2893 7046 2945 7098
rect 2957 7046 3009 7098
rect 3021 7046 3073 7098
rect 3085 7046 3137 7098
rect 3149 7046 3201 7098
rect 6780 7046 6832 7098
rect 6844 7046 6896 7098
rect 6908 7046 6960 7098
rect 6972 7046 7024 7098
rect 7036 7046 7088 7098
rect 10667 7046 10719 7098
rect 10731 7046 10783 7098
rect 10795 7046 10847 7098
rect 10859 7046 10911 7098
rect 10923 7046 10975 7098
rect 14554 7046 14606 7098
rect 14618 7046 14670 7098
rect 14682 7046 14734 7098
rect 14746 7046 14798 7098
rect 14810 7046 14862 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 2596 6944 2648 6996
rect 2780 6944 2832 6996
rect 3424 6944 3476 6996
rect 11060 6987 11112 6996
rect 11060 6953 11069 6987
rect 11069 6953 11103 6987
rect 11103 6953 11112 6987
rect 11060 6944 11112 6953
rect 14004 6944 14056 6996
rect 5356 6876 5408 6928
rect 5908 6876 5960 6928
rect 2596 6672 2648 6724
rect 2872 6740 2924 6792
rect 3424 6808 3476 6860
rect 5172 6808 5224 6860
rect 5264 6740 5316 6792
rect 11244 6876 11296 6928
rect 11888 6876 11940 6928
rect 12164 6876 12216 6928
rect 7380 6851 7432 6860
rect 7380 6817 7389 6851
rect 7389 6817 7423 6851
rect 7423 6817 7432 6851
rect 7380 6808 7432 6817
rect 9864 6740 9916 6792
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 6552 6672 6604 6724
rect 11244 6740 11296 6792
rect 4528 6604 4580 6656
rect 6368 6604 6420 6656
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 7564 6604 7616 6656
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 11428 6672 11480 6724
rect 11980 6808 12032 6860
rect 12348 6808 12400 6860
rect 13912 6851 13964 6860
rect 13912 6817 13921 6851
rect 13921 6817 13955 6851
rect 13955 6817 13964 6851
rect 13912 6808 13964 6817
rect 14280 6672 14332 6724
rect 15384 6672 15436 6724
rect 11152 6604 11204 6656
rect 11796 6604 11848 6656
rect 15844 6647 15896 6656
rect 15844 6613 15853 6647
rect 15853 6613 15887 6647
rect 15887 6613 15896 6647
rect 15844 6604 15896 6613
rect 4836 6502 4888 6554
rect 4900 6502 4952 6554
rect 4964 6502 5016 6554
rect 5028 6502 5080 6554
rect 5092 6502 5144 6554
rect 8723 6502 8775 6554
rect 8787 6502 8839 6554
rect 8851 6502 8903 6554
rect 8915 6502 8967 6554
rect 8979 6502 9031 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 16497 6502 16549 6554
rect 16561 6502 16613 6554
rect 16625 6502 16677 6554
rect 16689 6502 16741 6554
rect 16753 6502 16805 6554
rect 6920 6400 6972 6452
rect 7288 6400 7340 6452
rect 4528 6332 4580 6384
rect 5264 6332 5316 6384
rect 7104 6332 7156 6384
rect 9496 6332 9548 6384
rect 15844 6400 15896 6452
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 11336 6264 11388 6316
rect 11796 6264 11848 6316
rect 4528 6239 4580 6248
rect 4528 6205 4537 6239
rect 4537 6205 4571 6239
rect 4571 6205 4580 6239
rect 4528 6196 4580 6205
rect 5724 6196 5776 6248
rect 6644 6239 6696 6248
rect 6644 6205 6653 6239
rect 6653 6205 6687 6239
rect 6687 6205 6696 6239
rect 6644 6196 6696 6205
rect 3240 6103 3292 6112
rect 3240 6069 3249 6103
rect 3249 6069 3283 6103
rect 3283 6069 3292 6103
rect 3240 6060 3292 6069
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 12164 6264 12216 6316
rect 12256 6264 12308 6316
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 14924 6239 14976 6248
rect 14924 6205 14933 6239
rect 14933 6205 14967 6239
rect 14967 6205 14976 6239
rect 14924 6196 14976 6205
rect 14280 6103 14332 6112
rect 14280 6069 14289 6103
rect 14289 6069 14323 6103
rect 14323 6069 14332 6103
rect 14280 6060 14332 6069
rect 2893 5958 2945 6010
rect 2957 5958 3009 6010
rect 3021 5958 3073 6010
rect 3085 5958 3137 6010
rect 3149 5958 3201 6010
rect 6780 5958 6832 6010
rect 6844 5958 6896 6010
rect 6908 5958 6960 6010
rect 6972 5958 7024 6010
rect 7036 5958 7088 6010
rect 10667 5958 10719 6010
rect 10731 5958 10783 6010
rect 10795 5958 10847 6010
rect 10859 5958 10911 6010
rect 10923 5958 10975 6010
rect 14554 5958 14606 6010
rect 14618 5958 14670 6010
rect 14682 5958 14734 6010
rect 14746 5958 14798 6010
rect 14810 5958 14862 6010
rect 2964 5856 3016 5908
rect 3424 5856 3476 5908
rect 4528 5856 4580 5908
rect 5264 5856 5316 5908
rect 6644 5856 6696 5908
rect 7104 5856 7156 5908
rect 8668 5856 8720 5908
rect 8852 5856 8904 5908
rect 9312 5856 9364 5908
rect 6460 5788 6512 5840
rect 3332 5720 3384 5772
rect 2780 5652 2832 5704
rect 4436 5652 4488 5704
rect 5172 5652 5224 5704
rect 5448 5720 5500 5772
rect 9496 5720 9548 5772
rect 12256 5856 12308 5908
rect 12072 5788 12124 5840
rect 11428 5720 11480 5772
rect 14280 5856 14332 5908
rect 16120 5899 16172 5908
rect 16120 5865 16129 5899
rect 16129 5865 16163 5899
rect 16163 5865 16172 5899
rect 16120 5856 16172 5865
rect 4068 5584 4120 5636
rect 12624 5652 12676 5704
rect 13636 5652 13688 5704
rect 7564 5584 7616 5636
rect 8300 5584 8352 5636
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 3976 5559 4028 5568
rect 3976 5525 3985 5559
rect 3985 5525 4019 5559
rect 4019 5525 4028 5559
rect 3976 5516 4028 5525
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 10416 5627 10468 5636
rect 10416 5593 10425 5627
rect 10425 5593 10459 5627
rect 10459 5593 10468 5627
rect 10416 5584 10468 5593
rect 16948 5584 17000 5636
rect 11980 5559 12032 5568
rect 11980 5525 11989 5559
rect 11989 5525 12023 5559
rect 12023 5525 12032 5559
rect 11980 5516 12032 5525
rect 12348 5559 12400 5568
rect 12348 5525 12357 5559
rect 12357 5525 12391 5559
rect 12391 5525 12400 5559
rect 12348 5516 12400 5525
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 4836 5414 4888 5466
rect 4900 5414 4952 5466
rect 4964 5414 5016 5466
rect 5028 5414 5080 5466
rect 5092 5414 5144 5466
rect 8723 5414 8775 5466
rect 8787 5414 8839 5466
rect 8851 5414 8903 5466
rect 8915 5414 8967 5466
rect 8979 5414 9031 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 16497 5414 16549 5466
rect 16561 5414 16613 5466
rect 16625 5414 16677 5466
rect 16689 5414 16741 5466
rect 16753 5414 16805 5466
rect 3056 5312 3108 5364
rect 8300 5312 8352 5364
rect 9588 5312 9640 5364
rect 10416 5312 10468 5364
rect 11980 5312 12032 5364
rect 2504 5244 2556 5296
rect 3240 5244 3292 5296
rect 3976 5244 4028 5296
rect 4712 5176 4764 5228
rect 9496 5244 9548 5296
rect 2412 5108 2464 5160
rect 2596 5108 2648 5160
rect 9772 5176 9824 5228
rect 12072 5244 12124 5296
rect 11612 5219 11664 5228
rect 11612 5185 11621 5219
rect 11621 5185 11655 5219
rect 11655 5185 11664 5219
rect 11612 5176 11664 5185
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 1676 4972 1728 5024
rect 4160 4972 4212 5024
rect 5264 5015 5316 5024
rect 5264 4981 5273 5015
rect 5273 4981 5307 5015
rect 5307 4981 5316 5015
rect 5264 4972 5316 4981
rect 7380 4972 7432 5024
rect 12164 5176 12216 5228
rect 14372 5244 14424 5296
rect 13912 5176 13964 5228
rect 15752 5176 15804 5228
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 15936 5015 15988 5024
rect 15936 4981 15945 5015
rect 15945 4981 15979 5015
rect 15979 4981 15988 5015
rect 15936 4972 15988 4981
rect 2893 4870 2945 4922
rect 2957 4870 3009 4922
rect 3021 4870 3073 4922
rect 3085 4870 3137 4922
rect 3149 4870 3201 4922
rect 6780 4870 6832 4922
rect 6844 4870 6896 4922
rect 6908 4870 6960 4922
rect 6972 4870 7024 4922
rect 7036 4870 7088 4922
rect 10667 4870 10719 4922
rect 10731 4870 10783 4922
rect 10795 4870 10847 4922
rect 10859 4870 10911 4922
rect 10923 4870 10975 4922
rect 14554 4870 14606 4922
rect 14618 4870 14670 4922
rect 14682 4870 14734 4922
rect 14746 4870 14798 4922
rect 14810 4870 14862 4922
rect 4712 4811 4764 4820
rect 4712 4777 4721 4811
rect 4721 4777 4755 4811
rect 4755 4777 4764 4811
rect 4712 4768 4764 4777
rect 5264 4768 5316 4820
rect 5448 4768 5500 4820
rect 7380 4768 7432 4820
rect 9772 4811 9824 4820
rect 9772 4777 9781 4811
rect 9781 4777 9815 4811
rect 9815 4777 9824 4811
rect 9772 4768 9824 4777
rect 13636 4768 13688 4820
rect 15936 4768 15988 4820
rect 2504 4700 2556 4752
rect 1676 4607 1728 4616
rect 1676 4573 1710 4607
rect 1710 4573 1728 4607
rect 1676 4564 1728 4573
rect 2412 4564 2464 4616
rect 5356 4675 5408 4684
rect 5356 4641 5365 4675
rect 5365 4641 5399 4675
rect 5399 4641 5408 4675
rect 5356 4632 5408 4641
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4436 4564 4488 4616
rect 5172 4564 5224 4616
rect 13820 4700 13872 4752
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 14924 4632 14976 4684
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 11796 4564 11848 4616
rect 12164 4564 12216 4616
rect 6460 4428 6512 4480
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 7748 4471 7800 4480
rect 7748 4437 7757 4471
rect 7757 4437 7791 4471
rect 7791 4437 7800 4471
rect 7748 4428 7800 4437
rect 9588 4428 9640 4480
rect 10140 4471 10192 4480
rect 10140 4437 10149 4471
rect 10149 4437 10183 4471
rect 10183 4437 10192 4471
rect 10140 4428 10192 4437
rect 14004 4428 14056 4480
rect 4836 4326 4888 4378
rect 4900 4326 4952 4378
rect 4964 4326 5016 4378
rect 5028 4326 5080 4378
rect 5092 4326 5144 4378
rect 8723 4326 8775 4378
rect 8787 4326 8839 4378
rect 8851 4326 8903 4378
rect 8915 4326 8967 4378
rect 8979 4326 9031 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 16497 4326 16549 4378
rect 16561 4326 16613 4378
rect 16625 4326 16677 4378
rect 16689 4326 16741 4378
rect 16753 4326 16805 4378
rect 5172 4267 5224 4276
rect 5172 4233 5181 4267
rect 5181 4233 5215 4267
rect 5215 4233 5224 4267
rect 5172 4224 5224 4233
rect 940 4156 992 4208
rect 3792 4156 3844 4208
rect 4436 4156 4488 4208
rect 7748 4156 7800 4208
rect 10140 4156 10192 4208
rect 2780 4088 2832 4140
rect 2412 4020 2464 4072
rect 6460 4088 6512 4140
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 5724 4020 5776 4029
rect 4436 3884 4488 3936
rect 5356 3952 5408 4004
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 12256 4088 12308 4140
rect 12348 4088 12400 4140
rect 13912 4156 13964 4208
rect 11060 3952 11112 4004
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 5264 3927 5316 3936
rect 5264 3893 5273 3927
rect 5273 3893 5307 3927
rect 5307 3893 5316 3927
rect 5264 3884 5316 3893
rect 12256 3884 12308 3936
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 15752 4020 15804 4072
rect 13728 3952 13780 4004
rect 2893 3782 2945 3834
rect 2957 3782 3009 3834
rect 3021 3782 3073 3834
rect 3085 3782 3137 3834
rect 3149 3782 3201 3834
rect 6780 3782 6832 3834
rect 6844 3782 6896 3834
rect 6908 3782 6960 3834
rect 6972 3782 7024 3834
rect 7036 3782 7088 3834
rect 10667 3782 10719 3834
rect 10731 3782 10783 3834
rect 10795 3782 10847 3834
rect 10859 3782 10911 3834
rect 10923 3782 10975 3834
rect 14554 3782 14606 3834
rect 14618 3782 14670 3834
rect 14682 3782 14734 3834
rect 14746 3782 14798 3834
rect 14810 3782 14862 3834
rect 3976 3680 4028 3732
rect 6644 3680 6696 3732
rect 10324 3723 10376 3732
rect 10324 3689 10333 3723
rect 10333 3689 10367 3723
rect 10367 3689 10376 3723
rect 10324 3680 10376 3689
rect 11060 3680 11112 3732
rect 11520 3680 11572 3732
rect 12532 3680 12584 3732
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 11888 3587 11940 3596
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 12256 3544 12308 3596
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4712 3476 4764 3528
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 4068 3408 4120 3460
rect 7288 3476 7340 3528
rect 13912 3680 13964 3732
rect 14188 3612 14240 3664
rect 8300 3408 8352 3460
rect 8576 3408 8628 3460
rect 2780 3383 2832 3392
rect 2780 3349 2789 3383
rect 2789 3349 2823 3383
rect 2823 3349 2832 3383
rect 2780 3340 2832 3349
rect 3792 3340 3844 3392
rect 4712 3383 4764 3392
rect 4712 3349 4721 3383
rect 4721 3349 4755 3383
rect 4755 3349 4764 3383
rect 4712 3340 4764 3349
rect 5448 3383 5500 3392
rect 5448 3349 5457 3383
rect 5457 3349 5491 3383
rect 5491 3349 5500 3383
rect 5448 3340 5500 3349
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 10784 3383 10836 3392
rect 10784 3349 10793 3383
rect 10793 3349 10827 3383
rect 10827 3349 10836 3383
rect 10784 3340 10836 3349
rect 16120 3408 16172 3460
rect 4836 3238 4888 3290
rect 4900 3238 4952 3290
rect 4964 3238 5016 3290
rect 5028 3238 5080 3290
rect 5092 3238 5144 3290
rect 8723 3238 8775 3290
rect 8787 3238 8839 3290
rect 8851 3238 8903 3290
rect 8915 3238 8967 3290
rect 8979 3238 9031 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 16497 3238 16549 3290
rect 16561 3238 16613 3290
rect 16625 3238 16677 3290
rect 16689 3238 16741 3290
rect 16753 3238 16805 3290
rect 2780 3136 2832 3188
rect 3792 3179 3844 3188
rect 3792 3145 3801 3179
rect 3801 3145 3835 3179
rect 3835 3145 3844 3179
rect 3792 3136 3844 3145
rect 4068 3136 4120 3188
rect 5724 3136 5776 3188
rect 7472 3136 7524 3188
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 4712 3111 4764 3120
rect 4712 3077 4735 3111
rect 4735 3077 4764 3111
rect 4712 3068 4764 3077
rect 6460 3043 6512 3052
rect 6460 3009 6469 3043
rect 6469 3009 6503 3043
rect 6503 3009 6512 3043
rect 6460 3000 6512 3009
rect 7104 3000 7156 3052
rect 8300 3000 8352 3052
rect 8484 2975 8536 2984
rect 8484 2941 8493 2975
rect 8493 2941 8527 2975
rect 8527 2941 8536 2975
rect 8484 2932 8536 2941
rect 11704 3136 11756 3188
rect 13176 3136 13228 3188
rect 9588 3068 9640 3120
rect 10508 3000 10560 3052
rect 11888 3000 11940 3052
rect 12256 3043 12308 3052
rect 12256 3009 12290 3043
rect 12290 3009 12308 3043
rect 12256 3000 12308 3009
rect 4252 2839 4304 2848
rect 4252 2805 4261 2839
rect 4261 2805 4295 2839
rect 4295 2805 4304 2839
rect 4252 2796 4304 2805
rect 7932 2839 7984 2848
rect 7932 2805 7941 2839
rect 7941 2805 7975 2839
rect 7975 2805 7984 2839
rect 7932 2796 7984 2805
rect 10416 2796 10468 2848
rect 10784 2796 10836 2848
rect 2893 2694 2945 2746
rect 2957 2694 3009 2746
rect 3021 2694 3073 2746
rect 3085 2694 3137 2746
rect 3149 2694 3201 2746
rect 6780 2694 6832 2746
rect 6844 2694 6896 2746
rect 6908 2694 6960 2746
rect 6972 2694 7024 2746
rect 7036 2694 7088 2746
rect 10667 2694 10719 2746
rect 10731 2694 10783 2746
rect 10795 2694 10847 2746
rect 10859 2694 10911 2746
rect 10923 2694 10975 2746
rect 14554 2694 14606 2746
rect 14618 2694 14670 2746
rect 14682 2694 14734 2746
rect 14746 2694 14798 2746
rect 14810 2694 14862 2746
rect 2780 2592 2832 2644
rect 3884 2592 3936 2644
rect 4712 2592 4764 2644
rect 6368 2592 6420 2644
rect 7104 2592 7156 2644
rect 7932 2592 7984 2644
rect 8392 2592 8444 2644
rect 10508 2635 10560 2644
rect 10508 2601 10517 2635
rect 10517 2601 10551 2635
rect 10551 2601 10560 2635
rect 10508 2592 10560 2601
rect 12256 2592 12308 2644
rect 12440 2592 12492 2644
rect 16120 2635 16172 2644
rect 16120 2601 16129 2635
rect 16129 2601 16163 2635
rect 16163 2601 16172 2635
rect 16120 2592 16172 2601
rect 2596 2456 2648 2508
rect 4252 2456 4304 2508
rect 11704 2524 11756 2576
rect 20 2388 72 2440
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 5724 2388 5776 2440
rect 6460 2388 6512 2440
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 3792 2320 3844 2372
rect 4068 2363 4120 2372
rect 4068 2329 4077 2363
rect 4077 2329 4111 2363
rect 4111 2329 4120 2363
rect 4068 2320 4120 2329
rect 10048 2388 10100 2440
rect 11980 2456 12032 2508
rect 5172 2252 5224 2304
rect 10416 2320 10468 2372
rect 12164 2431 12216 2440
rect 12164 2397 12173 2431
rect 12173 2397 12207 2431
rect 12207 2397 12216 2431
rect 12164 2388 12216 2397
rect 11796 2252 11848 2304
rect 13360 2320 13412 2372
rect 15660 2363 15712 2372
rect 15660 2329 15669 2363
rect 15669 2329 15703 2363
rect 15703 2329 15712 2363
rect 15660 2320 15712 2329
rect 16396 2252 16448 2304
rect 4836 2150 4888 2202
rect 4900 2150 4952 2202
rect 4964 2150 5016 2202
rect 5028 2150 5080 2202
rect 5092 2150 5144 2202
rect 8723 2150 8775 2202
rect 8787 2150 8839 2202
rect 8851 2150 8903 2202
rect 8915 2150 8967 2202
rect 8979 2150 9031 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 16497 2150 16549 2202
rect 16561 2150 16613 2202
rect 16625 2150 16677 2202
rect 16689 2150 16741 2202
rect 16753 2150 16805 2202
<< metal2 >>
rect 18 19145 74 19945
rect 3882 19258 3938 19945
rect 3620 19230 3938 19258
rect 32 17338 60 19145
rect 20 17332 72 17338
rect 20 17274 72 17280
rect 3620 17270 3648 19230
rect 3882 19145 3938 19230
rect 7746 19145 7802 19945
rect 11610 19145 11666 19945
rect 15474 19145 15530 19945
rect 4836 17436 5144 17445
rect 4836 17434 4842 17436
rect 4898 17434 4922 17436
rect 4978 17434 5002 17436
rect 5058 17434 5082 17436
rect 5138 17434 5144 17436
rect 4898 17382 4900 17434
rect 5080 17382 5082 17434
rect 4836 17380 4842 17382
rect 4898 17380 4922 17382
rect 4978 17380 5002 17382
rect 5058 17380 5082 17382
rect 5138 17380 5144 17382
rect 4836 17371 5144 17380
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 3608 17264 3660 17270
rect 3608 17206 3660 17212
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 940 16584 992 16590
rect 940 16526 992 16532
rect 952 16425 980 16526
rect 938 16416 994 16425
rect 938 16351 994 16360
rect 1504 15162 1532 17138
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 2893 16892 3201 16901
rect 2893 16890 2899 16892
rect 2955 16890 2979 16892
rect 3035 16890 3059 16892
rect 3115 16890 3139 16892
rect 3195 16890 3201 16892
rect 2955 16838 2957 16890
rect 3137 16838 3139 16890
rect 2893 16836 2899 16838
rect 2955 16836 2979 16838
rect 3035 16836 3059 16838
rect 3115 16836 3139 16838
rect 3195 16836 3201 16838
rect 2893 16827 3201 16836
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 2148 16250 2176 16458
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2700 16250 2728 16390
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2792 16114 2820 16390
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 14482 1440 14894
rect 1688 14618 1716 14962
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 2332 14414 2360 15098
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12345 1624 12582
rect 1582 12336 1638 12345
rect 1780 12306 1808 14010
rect 2608 13938 2636 14214
rect 2792 14074 2820 16050
rect 2893 15804 3201 15813
rect 2893 15802 2899 15804
rect 2955 15802 2979 15804
rect 3035 15802 3059 15804
rect 3115 15802 3139 15804
rect 3195 15802 3201 15804
rect 2955 15750 2957 15802
rect 3137 15750 3139 15802
rect 2893 15748 2899 15750
rect 2955 15748 2979 15750
rect 3035 15748 3059 15750
rect 3115 15748 3139 15750
rect 3195 15748 3201 15750
rect 2893 15739 3201 15748
rect 2893 14716 3201 14725
rect 2893 14714 2899 14716
rect 2955 14714 2979 14716
rect 3035 14714 3059 14716
rect 3115 14714 3139 14716
rect 3195 14714 3201 14716
rect 2955 14662 2957 14714
rect 3137 14662 3139 14714
rect 2893 14660 2899 14662
rect 2955 14660 2979 14662
rect 3035 14660 3059 14662
rect 3115 14660 3139 14662
rect 3195 14660 3201 14662
rect 2893 14651 3201 14660
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3160 14074 3188 14350
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2893 13628 3201 13637
rect 2893 13626 2899 13628
rect 2955 13626 2979 13628
rect 3035 13626 3059 13628
rect 3115 13626 3139 13628
rect 3195 13626 3201 13628
rect 2955 13574 2957 13626
rect 3137 13574 3139 13626
rect 2893 13572 2899 13574
rect 2955 13572 2979 13574
rect 3035 13572 3059 13574
rect 3115 13572 3139 13574
rect 3195 13572 3201 13574
rect 2893 13563 3201 13572
rect 3252 13410 3280 16730
rect 3344 14414 3372 16934
rect 3804 16726 3832 17070
rect 3896 16794 3924 17138
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3436 15706 3464 15982
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3712 15502 3740 16050
rect 3804 16046 3832 16662
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4172 16046 4200 16594
rect 4632 16590 4660 17274
rect 7760 17270 7788 19145
rect 8723 17436 9031 17445
rect 8723 17434 8729 17436
rect 8785 17434 8809 17436
rect 8865 17434 8889 17436
rect 8945 17434 8969 17436
rect 9025 17434 9031 17436
rect 8785 17382 8787 17434
rect 8967 17382 8969 17434
rect 8723 17380 8729 17382
rect 8785 17380 8809 17382
rect 8865 17380 8889 17382
rect 8945 17380 8969 17382
rect 9025 17380 9031 17382
rect 8723 17371 9031 17380
rect 11624 17270 11652 19145
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12610 17371 12918 17380
rect 15488 17338 15516 19145
rect 15934 17776 15990 17785
rect 15934 17711 15990 17720
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15948 17270 15976 17711
rect 16497 17436 16805 17445
rect 16497 17434 16503 17436
rect 16559 17434 16583 17436
rect 16639 17434 16663 17436
rect 16719 17434 16743 17436
rect 16799 17434 16805 17436
rect 16559 17382 16561 17434
rect 16741 17382 16743 17434
rect 16497 17380 16503 17382
rect 16559 17380 16583 17382
rect 16639 17380 16663 17382
rect 16719 17380 16743 17382
rect 16799 17380 16805 17382
rect 16497 17371 16805 17380
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 4836 16348 5144 16357
rect 4836 16346 4842 16348
rect 4898 16346 4922 16348
rect 4978 16346 5002 16348
rect 5058 16346 5082 16348
rect 5138 16346 5144 16348
rect 4898 16294 4900 16346
rect 5080 16294 5082 16346
rect 4836 16292 4842 16294
rect 4898 16292 4922 16294
rect 4978 16292 5002 16294
rect 5058 16292 5082 16294
rect 5138 16292 5144 16294
rect 4836 16283 5144 16292
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3712 14414 3740 15438
rect 3804 14482 3832 15982
rect 4172 15314 4200 15982
rect 4724 15706 4752 15982
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 5184 15638 5212 16390
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 5276 15502 5304 16934
rect 6780 16892 7088 16901
rect 6780 16890 6786 16892
rect 6842 16890 6866 16892
rect 6922 16890 6946 16892
rect 7002 16890 7026 16892
rect 7082 16890 7088 16892
rect 6842 16838 6844 16890
rect 7024 16838 7026 16890
rect 6780 16836 6786 16838
rect 6842 16836 6866 16838
rect 6922 16836 6946 16838
rect 7002 16836 7026 16838
rect 7082 16836 7088 16838
rect 6780 16827 7088 16836
rect 7116 16794 7144 17138
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6472 16250 6500 16594
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 6748 16250 6776 16458
rect 7300 16250 7328 16458
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 4908 15366 4936 15438
rect 4080 15286 4200 15314
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3332 14408 3384 14414
rect 3700 14408 3752 14414
rect 3384 14368 3464 14396
rect 3332 14350 3384 14356
rect 3436 13870 3464 14368
rect 3700 14350 3752 14356
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3620 14074 3648 14214
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 2884 13382 3280 13410
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12850 2728 13126
rect 2884 12850 2912 13382
rect 3056 13184 3108 13190
rect 3332 13184 3384 13190
rect 3108 13144 3280 13172
rect 3056 13126 3108 13132
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 1582 12271 1638 12280
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11150 1900 11494
rect 2056 11150 2084 12378
rect 2332 12306 2360 12786
rect 2884 12730 2912 12786
rect 2700 12702 2912 12730
rect 2700 12374 2728 12702
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2792 12238 2820 12582
rect 2893 12540 3201 12549
rect 2893 12538 2899 12540
rect 2955 12538 2979 12540
rect 3035 12538 3059 12540
rect 3115 12538 3139 12540
rect 3195 12538 3201 12540
rect 2955 12486 2957 12538
rect 3137 12486 3139 12538
rect 2893 12484 2899 12486
rect 2955 12484 2979 12486
rect 3035 12484 3059 12486
rect 3115 12484 3139 12486
rect 3195 12484 3201 12486
rect 2893 12475 3201 12484
rect 3252 12442 3280 13144
rect 3332 13126 3384 13132
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11150 2268 11494
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1688 10742 1716 10950
rect 1676 10736 1728 10742
rect 1676 10678 1728 10684
rect 2056 10674 2084 11086
rect 2792 10810 2820 11698
rect 2893 11452 3201 11461
rect 2893 11450 2899 11452
rect 2955 11450 2979 11452
rect 3035 11450 3059 11452
rect 3115 11450 3139 11452
rect 3195 11450 3201 11452
rect 2955 11398 2957 11450
rect 3137 11398 3139 11450
rect 2893 11396 2899 11398
rect 2955 11396 2979 11398
rect 3035 11396 3059 11398
rect 3115 11396 3139 11398
rect 3195 11396 3201 11398
rect 2893 11387 3201 11396
rect 3344 11354 3372 13126
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3344 10810 3372 11290
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2056 10130 2084 10610
rect 2893 10364 3201 10373
rect 2893 10362 2899 10364
rect 2955 10362 2979 10364
rect 3035 10362 3059 10364
rect 3115 10362 3139 10364
rect 3195 10362 3201 10364
rect 2955 10310 2957 10362
rect 3137 10310 3139 10362
rect 2893 10308 2899 10310
rect 2955 10308 2979 10310
rect 3035 10308 3059 10310
rect 3115 10308 3139 10310
rect 3195 10308 3201 10310
rect 2893 10299 3201 10308
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1504 8566 1532 9522
rect 1688 9178 1716 9522
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2792 9178 2820 9386
rect 2893 9276 3201 9285
rect 2893 9274 2899 9276
rect 2955 9274 2979 9276
rect 3035 9274 3059 9276
rect 3115 9274 3139 9276
rect 3195 9274 3201 9276
rect 2955 9222 2957 9274
rect 3137 9222 3139 9274
rect 2893 9220 2899 9222
rect 2955 9220 2979 9222
rect 3035 9220 3059 9222
rect 3115 9220 3139 9222
rect 3195 9220 3201 9222
rect 2893 9211 3201 9220
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8634 2360 8774
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 1492 8560 1544 8566
rect 1492 8502 1544 8508
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1504 7410 1532 8502
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1688 7002 1716 7346
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 2516 6882 2544 8434
rect 2608 7954 2636 8978
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2792 8090 2820 8502
rect 2893 8188 3201 8197
rect 2893 8186 2899 8188
rect 2955 8186 2979 8188
rect 3035 8186 3059 8188
rect 3115 8186 3139 8188
rect 3195 8186 3201 8188
rect 2955 8134 2957 8186
rect 3137 8134 3139 8186
rect 2893 8132 2899 8134
rect 2955 8132 2979 8134
rect 3035 8132 3059 8134
rect 3115 8132 3139 8134
rect 3195 8132 3201 8134
rect 2893 8123 3201 8132
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2608 7002 2636 7890
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2792 7002 2820 7482
rect 3436 7426 3464 13806
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3528 10470 3556 12718
rect 3712 11150 3740 14350
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3896 13870 3924 14214
rect 4080 13870 4108 15286
rect 4836 15260 5144 15269
rect 4836 15258 4842 15260
rect 4898 15258 4922 15260
rect 4978 15258 5002 15260
rect 5058 15258 5082 15260
rect 5138 15258 5144 15260
rect 4898 15206 4900 15258
rect 5080 15206 5082 15258
rect 4836 15204 4842 15206
rect 4898 15204 4922 15206
rect 4978 15204 5002 15206
rect 5058 15204 5082 15206
rect 5138 15204 5144 15206
rect 4836 15195 5144 15204
rect 5172 14544 5224 14550
rect 5172 14486 5224 14492
rect 4896 14408 4948 14414
rect 4724 14368 4896 14396
rect 4724 14074 4752 14368
rect 4896 14350 4948 14356
rect 4836 14172 5144 14181
rect 4836 14170 4842 14172
rect 4898 14170 4922 14172
rect 4978 14170 5002 14172
rect 5058 14170 5082 14172
rect 5138 14170 5144 14172
rect 4898 14118 4900 14170
rect 5080 14118 5082 14170
rect 4836 14116 4842 14118
rect 4898 14116 4922 14118
rect 4978 14116 5002 14118
rect 5058 14116 5082 14118
rect 5138 14116 5144 14118
rect 4836 14107 5144 14116
rect 5184 14074 5212 14486
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11558 3924 12174
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3712 10674 3740 11086
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3620 9722 3648 9998
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3344 7398 3464 7426
rect 2893 7100 3201 7109
rect 2893 7098 2899 7100
rect 2955 7098 2979 7100
rect 3035 7098 3059 7100
rect 3115 7098 3139 7100
rect 3195 7098 3201 7100
rect 2955 7046 2957 7098
rect 3137 7046 3139 7098
rect 2893 7044 2899 7046
rect 2955 7044 2979 7046
rect 3035 7044 3059 7046
rect 3115 7044 3139 7046
rect 3195 7044 3201 7046
rect 2893 7035 3201 7044
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2516 6854 2820 6882
rect 2792 6746 2820 6854
rect 2872 6792 2924 6798
rect 2792 6740 2872 6746
rect 2792 6734 2924 6740
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2792 6718 2912 6734
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4622 1716 4966
rect 2424 4622 2452 5102
rect 2516 4758 2544 5238
rect 2608 5166 2636 6666
rect 2792 5710 2820 6718
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 2893 6012 3201 6021
rect 2893 6010 2899 6012
rect 2955 6010 2979 6012
rect 3035 6010 3059 6012
rect 3115 6010 3139 6012
rect 3195 6010 3201 6012
rect 2955 5958 2957 6010
rect 3137 5958 3139 6010
rect 2893 5956 2899 5958
rect 2955 5956 2979 5958
rect 3035 5956 3059 5958
rect 3115 5956 3139 5958
rect 3195 5956 3201 5958
rect 2893 5947 3201 5956
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2976 5250 3004 5850
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 5370 3096 5510
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3252 5302 3280 6054
rect 3344 5778 3372 7398
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3804 7290 3832 11154
rect 3896 10674 3924 11494
rect 3988 11286 4016 11834
rect 4080 11354 4108 13806
rect 4724 13394 4752 13874
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5276 13530 5304 13806
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4724 12986 4752 13330
rect 4836 13084 5144 13093
rect 4836 13082 4842 13084
rect 4898 13082 4922 13084
rect 4978 13082 5002 13084
rect 5058 13082 5082 13084
rect 5138 13082 5144 13084
rect 4898 13030 4900 13082
rect 5080 13030 5082 13082
rect 4836 13028 4842 13030
rect 4898 13028 4922 13030
rect 4978 13028 5002 13030
rect 5058 13028 5082 13030
rect 5138 13028 5144 13030
rect 4836 13019 5144 13028
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4172 12442 4200 12854
rect 5368 12442 5396 13874
rect 5460 12753 5488 15302
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5644 13938 5672 14350
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5644 13394 5672 13670
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5446 12744 5502 12753
rect 5446 12679 5502 12688
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 4836 11996 5144 12005
rect 4836 11994 4842 11996
rect 4898 11994 4922 11996
rect 4978 11994 5002 11996
rect 5058 11994 5082 11996
rect 5138 11994 5144 11996
rect 4898 11942 4900 11994
rect 5080 11942 5082 11994
rect 4836 11940 4842 11942
rect 4898 11940 4922 11942
rect 4978 11940 5002 11942
rect 5058 11940 5082 11942
rect 5138 11940 5144 11942
rect 4836 11931 5144 11940
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4080 10470 4108 11290
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4172 10810 4200 10950
rect 4724 10810 4752 11018
rect 4836 10908 5144 10917
rect 4836 10906 4842 10908
rect 4898 10906 4922 10908
rect 4978 10906 5002 10908
rect 5058 10906 5082 10908
rect 5138 10906 5144 10908
rect 4898 10854 4900 10906
rect 5080 10854 5082 10906
rect 4836 10852 4842 10854
rect 4898 10852 4922 10854
rect 4978 10852 5002 10854
rect 5058 10852 5082 10854
rect 5138 10852 5144 10854
rect 4836 10843 5144 10852
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4356 9654 4384 10542
rect 5368 10198 5396 10542
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4540 9722 4568 9930
rect 4836 9820 5144 9829
rect 4836 9818 4842 9820
rect 4898 9818 4922 9820
rect 4978 9818 5002 9820
rect 5058 9818 5082 9820
rect 5138 9818 5144 9820
rect 4898 9766 4900 9818
rect 5080 9766 5082 9818
rect 4836 9764 4842 9766
rect 4898 9764 4922 9766
rect 4978 9764 5002 9766
rect 5058 9764 5082 9766
rect 5138 9764 5144 9766
rect 4836 9755 5144 9764
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3896 8634 3924 9522
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3988 8498 4016 8774
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 4172 7954 4200 9454
rect 4356 9042 4384 9590
rect 5368 9058 5396 10134
rect 4344 9036 4396 9042
rect 5276 9030 5396 9058
rect 5460 9042 5488 12679
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5552 10266 5580 12242
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5644 10062 5672 13330
rect 6196 13326 6224 15846
rect 6288 15706 6316 16118
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 6780 15804 7088 15813
rect 6780 15802 6786 15804
rect 6842 15802 6866 15804
rect 6922 15802 6946 15804
rect 7002 15802 7026 15804
rect 7082 15802 7088 15804
rect 6842 15750 6844 15802
rect 7024 15750 7026 15802
rect 6780 15748 6786 15750
rect 6842 15748 6866 15750
rect 6922 15748 6946 15750
rect 7002 15748 7026 15750
rect 7082 15748 7088 15750
rect 6780 15739 7088 15748
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 7668 15162 7696 16050
rect 7944 15502 7972 16050
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 6780 14716 7088 14725
rect 6780 14714 6786 14716
rect 6842 14714 6866 14716
rect 6922 14714 6946 14716
rect 7002 14714 7026 14716
rect 7082 14714 7088 14716
rect 6842 14662 6844 14714
rect 7024 14662 7026 14714
rect 6780 14660 6786 14662
rect 6842 14660 6866 14662
rect 6922 14660 6946 14662
rect 7002 14660 7026 14662
rect 7082 14660 7088 14662
rect 6780 14651 7088 14660
rect 7484 13938 7512 14758
rect 7760 14618 7788 14962
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7944 14414 7972 15438
rect 8036 15366 8064 16934
rect 8128 16250 8156 16934
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 8312 15162 8340 17002
rect 9324 16794 9352 17138
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8404 16250 8432 16526
rect 9416 16454 9444 17070
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 8723 16348 9031 16357
rect 8723 16346 8729 16348
rect 8785 16346 8809 16348
rect 8865 16346 8889 16348
rect 8945 16346 8969 16348
rect 9025 16346 9031 16348
rect 8785 16294 8787 16346
rect 8967 16294 8969 16346
rect 8723 16292 8729 16294
rect 8785 16292 8809 16294
rect 8865 16292 8889 16294
rect 8945 16292 8969 16294
rect 9025 16292 9031 16294
rect 8723 16283 9031 16292
rect 9416 16250 9444 16390
rect 9784 16250 9812 16458
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 6780 13628 7088 13637
rect 6780 13626 6786 13628
rect 6842 13626 6866 13628
rect 6922 13626 6946 13628
rect 7002 13626 7026 13628
rect 7082 13626 7088 13628
rect 6842 13574 6844 13626
rect 7024 13574 7026 13626
rect 6780 13572 6786 13574
rect 6842 13572 6866 13574
rect 6922 13572 6946 13574
rect 7002 13572 7026 13574
rect 7082 13572 7088 13574
rect 6780 13563 7088 13572
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 6196 12986 6224 13262
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 12220 5764 12582
rect 5920 12434 5948 12718
rect 5920 12406 6040 12434
rect 5908 12232 5960 12238
rect 5736 12192 5908 12220
rect 5908 12174 5960 12180
rect 6012 11354 6040 12406
rect 6380 11762 6408 12718
rect 6656 12442 6684 12718
rect 6780 12540 7088 12549
rect 6780 12538 6786 12540
rect 6842 12538 6866 12540
rect 6922 12538 6946 12540
rect 7002 12538 7026 12540
rect 7082 12538 7088 12540
rect 6842 12486 6844 12538
rect 7024 12486 7026 12538
rect 6780 12484 6786 12486
rect 6842 12484 6866 12486
rect 6922 12484 6946 12486
rect 7002 12484 7026 12486
rect 7082 12484 7088 12486
rect 6780 12475 7088 12484
rect 7116 12442 7144 12854
rect 7300 12442 7328 13262
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7668 12238 7696 14350
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7852 14074 7880 14214
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 8312 12986 8340 14486
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7944 12306 7972 12718
rect 8404 12646 8432 15846
rect 9416 15706 9444 15982
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 8723 15260 9031 15269
rect 8723 15258 8729 15260
rect 8785 15258 8809 15260
rect 8865 15258 8889 15260
rect 8945 15258 8969 15260
rect 9025 15258 9031 15260
rect 8785 15206 8787 15258
rect 8967 15206 8969 15258
rect 8723 15204 8729 15206
rect 8785 15204 8809 15206
rect 8865 15204 8889 15206
rect 8945 15204 8969 15206
rect 9025 15204 9031 15206
rect 8723 15195 9031 15204
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8588 14346 8616 14826
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8588 14074 8616 14282
rect 8723 14172 9031 14181
rect 8723 14170 8729 14172
rect 8785 14170 8809 14172
rect 8865 14170 8889 14172
rect 8945 14170 8969 14172
rect 9025 14170 9031 14172
rect 8785 14118 8787 14170
rect 8967 14118 8969 14170
rect 8723 14116 8729 14118
rect 8785 14116 8809 14118
rect 8865 14116 8889 14118
rect 8945 14116 8969 14118
rect 9025 14116 9031 14118
rect 8723 14107 9031 14116
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 9140 13802 9168 15030
rect 9232 13870 9260 15302
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 8723 13084 9031 13093
rect 8723 13082 8729 13084
rect 8785 13082 8809 13084
rect 8865 13082 8889 13084
rect 8945 13082 8969 13084
rect 9025 13082 9031 13084
rect 8785 13030 8787 13082
rect 8967 13030 8969 13082
rect 8723 13028 8729 13030
rect 8785 13028 8809 13030
rect 8865 13028 8889 13030
rect 8945 13028 8969 13030
rect 9025 13028 9031 13030
rect 8723 13019 9031 13028
rect 9140 12986 9168 13738
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8392 12640 8444 12646
rect 8588 12628 8616 12854
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8392 12582 8444 12588
rect 8496 12600 8616 12628
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 8128 12170 8156 12582
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6012 11150 6040 11290
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5828 10810 5856 11018
rect 6104 10810 6132 11222
rect 6380 11014 6408 11698
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6380 10130 6408 10950
rect 6656 10810 6684 11698
rect 7944 11558 7972 12038
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 6780 11452 7088 11461
rect 6780 11450 6786 11452
rect 6842 11450 6866 11452
rect 6922 11450 6946 11452
rect 7002 11450 7026 11452
rect 7082 11450 7088 11452
rect 6842 11398 6844 11450
rect 7024 11398 7026 11450
rect 6780 11396 6786 11398
rect 6842 11396 6866 11398
rect 6922 11396 6946 11398
rect 7002 11396 7026 11398
rect 7082 11396 7088 11398
rect 6780 11387 7088 11396
rect 7944 11150 7972 11494
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7024 10810 7052 10950
rect 7484 10810 7512 10950
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 6780 10364 7088 10373
rect 6780 10362 6786 10364
rect 6842 10362 6866 10364
rect 6922 10362 6946 10364
rect 7002 10362 7026 10364
rect 7082 10362 7088 10364
rect 6842 10310 6844 10362
rect 7024 10310 7026 10362
rect 6780 10308 6786 10310
rect 6842 10308 6866 10310
rect 6922 10308 6946 10310
rect 7002 10308 7026 10310
rect 7082 10308 7088 10310
rect 6780 10299 7088 10308
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6196 9654 6224 9862
rect 6380 9722 6408 10066
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6932 9722 6960 9930
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 5448 9036 5500 9042
rect 4396 8996 4476 9024
rect 4344 8978 4396 8984
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4080 7546 4108 7754
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 7546 4200 7686
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4448 7410 4476 8996
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 4836 8732 5144 8741
rect 4836 8730 4842 8732
rect 4898 8730 4922 8732
rect 4978 8730 5002 8732
rect 5058 8730 5082 8732
rect 5138 8730 5144 8732
rect 4898 8678 4900 8730
rect 5080 8678 5082 8730
rect 4836 8676 4842 8678
rect 4898 8676 4922 8678
rect 4978 8676 5002 8678
rect 5058 8676 5082 8678
rect 5138 8676 5144 8678
rect 4836 8667 5144 8676
rect 5184 8634 5212 8774
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 3436 7002 3464 7278
rect 3804 7262 3924 7290
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 5914 3464 6802
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 2792 5222 3004 5250
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 2596 5160 2648 5166
rect 2792 5114 2820 5222
rect 2596 5102 2648 5108
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 940 4208 992 4214
rect 938 4176 940 4185
rect 992 4176 994 4185
rect 938 4111 994 4120
rect 2424 4078 2452 4558
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2424 3058 2452 4014
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2608 2514 2636 5102
rect 2700 5086 2820 5114
rect 2700 4434 2728 5086
rect 2893 4924 3201 4933
rect 2893 4922 2899 4924
rect 2955 4922 2979 4924
rect 3035 4922 3059 4924
rect 3115 4922 3139 4924
rect 3195 4922 3201 4924
rect 2955 4870 2957 4922
rect 3137 4870 3139 4922
rect 2893 4868 2899 4870
rect 2955 4868 2979 4870
rect 3035 4868 3059 4870
rect 3115 4868 3139 4870
rect 3195 4868 3201 4870
rect 2893 4859 3201 4868
rect 3792 4480 3844 4486
rect 2700 4406 2820 4434
rect 3792 4422 3844 4428
rect 2792 4146 2820 4406
rect 3804 4214 3832 4422
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2893 3836 3201 3845
rect 2893 3834 2899 3836
rect 2955 3834 2979 3836
rect 3035 3834 3059 3836
rect 3115 3834 3139 3836
rect 3195 3834 3201 3836
rect 2955 3782 2957 3834
rect 3137 3782 3139 3834
rect 2893 3780 2899 3782
rect 2955 3780 2979 3782
rect 3035 3780 3059 3782
rect 3115 3780 3139 3782
rect 3195 3780 3201 3782
rect 2893 3771 3201 3780
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2792 3194 2820 3334
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2976 3074 3004 3470
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3804 3194 3832 3334
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 2792 3046 3004 3074
rect 2792 2650 2820 3046
rect 2893 2748 3201 2757
rect 2893 2746 2899 2748
rect 2955 2746 2979 2748
rect 3035 2746 3059 2748
rect 3115 2746 3139 2748
rect 3195 2746 3201 2748
rect 2955 2694 2957 2746
rect 3137 2694 3139 2746
rect 2893 2692 2899 2694
rect 2955 2692 2979 2694
rect 3035 2692 3059 2694
rect 3115 2692 3139 2694
rect 3195 2692 3201 2694
rect 2893 2683 3201 2692
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 32 800 60 2382
rect 3804 2378 3832 3130
rect 3896 3058 3924 7262
rect 4448 5710 4476 7346
rect 4540 7274 4568 8366
rect 4836 7644 5144 7653
rect 4836 7642 4842 7644
rect 4898 7642 4922 7644
rect 4978 7642 5002 7644
rect 5058 7642 5082 7644
rect 5138 7642 5144 7644
rect 4898 7590 4900 7642
rect 5080 7590 5082 7642
rect 4836 7588 4842 7590
rect 4898 7588 4922 7590
rect 4978 7588 5002 7590
rect 5058 7588 5082 7590
rect 5138 7588 5144 7590
rect 4836 7579 5144 7588
rect 5276 7290 5304 9030
rect 5448 8978 5500 8984
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5368 8090 5396 8910
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5828 7954 5856 8774
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 5184 7262 5304 7290
rect 4540 6662 4568 7210
rect 5184 6866 5212 7262
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5276 6798 5304 7142
rect 5368 6934 5396 7890
rect 6196 7886 6224 8230
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 5736 7546 5764 7822
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6390 4568 6598
rect 4836 6556 5144 6565
rect 4836 6554 4842 6556
rect 4898 6554 4922 6556
rect 4978 6554 5002 6556
rect 5058 6554 5082 6556
rect 5138 6554 5144 6556
rect 4898 6502 4900 6554
rect 5080 6502 5082 6554
rect 4836 6500 4842 6502
rect 4898 6500 4922 6502
rect 4978 6500 5002 6502
rect 5058 6500 5082 6502
rect 5138 6500 5144 6502
rect 4836 6491 5144 6500
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4540 5914 4568 6190
rect 5276 5914 5304 6326
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3988 5302 4016 5510
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3988 3738 4016 4558
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4080 3466 4108 5578
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 3534 4200 4966
rect 4448 4622 4476 5646
rect 4836 5468 5144 5477
rect 4836 5466 4842 5468
rect 4898 5466 4922 5468
rect 4978 5466 5002 5468
rect 5058 5466 5082 5468
rect 5138 5466 5144 5468
rect 4898 5414 4900 5466
rect 5080 5414 5082 5466
rect 4836 5412 4842 5414
rect 4898 5412 4922 5414
rect 4978 5412 5002 5414
rect 5058 5412 5082 5414
rect 5138 5412 5144 5414
rect 4836 5403 5144 5412
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4724 4826 4752 5170
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 5184 4706 5212 5646
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5276 4826 5304 4966
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5184 4678 5304 4706
rect 5368 4690 5396 6870
rect 5736 6254 5764 7346
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5920 6934 5948 7278
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6380 6322 6408 6598
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 6472 5846 6500 7822
rect 6564 6730 6592 9522
rect 6780 9276 7088 9285
rect 6780 9274 6786 9276
rect 6842 9274 6866 9276
rect 6922 9274 6946 9276
rect 7002 9274 7026 9276
rect 7082 9274 7088 9276
rect 6842 9222 6844 9274
rect 7024 9222 7026 9274
rect 6780 9220 6786 9222
rect 6842 9220 6866 9222
rect 6922 9220 6946 9222
rect 7002 9220 7026 9222
rect 7082 9220 7088 9222
rect 6780 9211 7088 9220
rect 7208 8566 7236 10542
rect 8036 9042 8064 11766
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8312 11370 8340 11494
rect 8220 11354 8340 11370
rect 8208 11348 8340 11354
rect 8260 11342 8340 11348
rect 8208 11290 8260 11296
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8312 10742 8340 11222
rect 8404 11098 8432 12582
rect 8496 12442 8524 12600
rect 8484 12436 8536 12442
rect 8680 12434 8708 12650
rect 8484 12378 8536 12384
rect 8588 12406 8708 12434
rect 8956 12434 8984 12786
rect 9232 12434 9260 13806
rect 9324 13394 9352 15030
rect 9600 14482 9628 15982
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9876 14618 9904 14894
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9416 14074 9444 14350
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9508 12986 9536 13194
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 8956 12406 9168 12434
rect 9232 12406 9536 12434
rect 8496 11218 8524 12378
rect 8588 11778 8616 12406
rect 8723 11996 9031 12005
rect 8723 11994 8729 11996
rect 8785 11994 8809 11996
rect 8865 11994 8889 11996
rect 8945 11994 8969 11996
rect 9025 11994 9031 11996
rect 8785 11942 8787 11994
rect 8967 11942 8969 11994
rect 8723 11940 8729 11942
rect 8785 11940 8809 11942
rect 8865 11940 8889 11942
rect 8945 11940 8969 11942
rect 9025 11940 9031 11942
rect 8723 11931 9031 11940
rect 9140 11778 9168 12406
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9324 11898 9352 12106
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 8588 11750 8708 11778
rect 9140 11750 9352 11778
rect 8680 11354 8708 11750
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9048 11234 9076 11290
rect 9220 11280 9272 11286
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8576 11212 8628 11218
rect 9048 11206 9168 11234
rect 9220 11222 9272 11228
rect 8576 11154 8628 11160
rect 8404 11070 8524 11098
rect 8496 11014 8524 11070
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10810 8524 10950
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8588 10606 8616 11154
rect 8723 10908 9031 10917
rect 8723 10906 8729 10908
rect 8785 10906 8809 10908
rect 8865 10906 8889 10908
rect 8945 10906 8969 10908
rect 9025 10906 9031 10908
rect 8785 10854 8787 10906
rect 8967 10854 8969 10906
rect 8723 10852 8729 10854
rect 8785 10852 8809 10854
rect 8865 10852 8889 10854
rect 8945 10852 8969 10854
rect 9025 10852 9031 10854
rect 8723 10843 9031 10852
rect 9140 10606 9168 11206
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 8128 9602 8156 10542
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8312 10266 8340 10474
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8128 9574 8248 9602
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8220 8974 8248 9574
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8312 9110 8340 9522
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7750 6684 8230
rect 6780 8188 7088 8197
rect 6780 8186 6786 8188
rect 6842 8186 6866 8188
rect 6922 8186 6946 8188
rect 7002 8186 7026 8188
rect 7082 8186 7088 8188
rect 6842 8134 6844 8186
rect 7024 8134 7026 8186
rect 6780 8132 6786 8134
rect 6842 8132 6866 8134
rect 6922 8132 6946 8134
rect 7002 8132 7026 8134
rect 7082 8132 7088 8134
rect 6780 8123 7088 8132
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 7116 7546 7144 8434
rect 8128 7886 8156 8774
rect 8220 8430 8248 8910
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 7392 7546 7420 7686
rect 8312 7546 8340 7686
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 6780 7100 7088 7109
rect 6780 7098 6786 7100
rect 6842 7098 6866 7100
rect 6922 7098 6946 7100
rect 7002 7098 7026 7100
rect 7082 7098 7088 7100
rect 6842 7046 6844 7098
rect 7024 7046 7026 7098
rect 6780 7044 6786 7046
rect 6842 7044 6866 7046
rect 6922 7044 6946 7046
rect 7002 7044 7026 7046
rect 7082 7044 7088 7046
rect 6780 7035 7088 7044
rect 7392 6866 7420 7482
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5460 4826 5488 5714
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4214 4476 4422
rect 4836 4380 5144 4389
rect 4836 4378 4842 4380
rect 4898 4378 4922 4380
rect 4978 4378 5002 4380
rect 5058 4378 5082 4380
rect 5138 4378 5144 4380
rect 4898 4326 4900 4378
rect 5080 4326 5082 4378
rect 4836 4324 4842 4326
rect 4898 4324 4922 4326
rect 4978 4324 5002 4326
rect 5058 4324 5082 4326
rect 5138 4324 5144 4326
rect 4836 4315 5144 4324
rect 5184 4282 5212 4558
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 5276 3942 5304 4678
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5368 4010 5396 4626
rect 6472 4486 6500 5782
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6472 4146 6500 4422
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 4448 3602 4476 3878
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4160 3528 4212 3534
rect 4712 3528 4764 3534
rect 4160 3470 4212 3476
rect 4632 3476 4712 3482
rect 4632 3470 4764 3476
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4632 3454 4752 3470
rect 4080 3194 4108 3402
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3896 2650 3924 2994
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 4264 2514 4292 2790
rect 4632 2774 4660 3454
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3126 4752 3334
rect 4836 3292 5144 3301
rect 4836 3290 4842 3292
rect 4898 3290 4922 3292
rect 4978 3290 5002 3292
rect 5058 3290 5082 3292
rect 5138 3290 5144 3292
rect 4898 3238 4900 3290
rect 5080 3238 5082 3290
rect 4836 3236 4842 3238
rect 4898 3236 4922 3238
rect 4978 3236 5002 3238
rect 5058 3236 5082 3238
rect 5138 3236 5144 3238
rect 4836 3227 5144 3236
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4632 2746 4752 2774
rect 4724 2650 4752 2746
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4080 1170 4108 2314
rect 5184 2310 5212 3470
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 2774 5488 3334
rect 5736 3194 5764 4014
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5368 2746 5488 2774
rect 5368 2446 5396 2746
rect 5736 2446 5764 3130
rect 6472 3058 6500 4082
rect 6460 3052 6512 3058
rect 6380 3012 6460 3040
rect 6380 2650 6408 3012
rect 6460 2994 6512 3000
rect 6564 2774 6592 6666
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 6932 6458 6960 6598
rect 7300 6458 7328 6598
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6656 5914 6684 6190
rect 6780 6012 7088 6021
rect 6780 6010 6786 6012
rect 6842 6010 6866 6012
rect 6922 6010 6946 6012
rect 7002 6010 7026 6012
rect 7082 6010 7088 6012
rect 6842 5958 6844 6010
rect 7024 5958 7026 6010
rect 6780 5956 6786 5958
rect 6842 5956 6866 5958
rect 6922 5956 6946 5958
rect 7002 5956 7026 5958
rect 7082 5956 7088 5958
rect 6780 5947 7088 5956
rect 7116 5914 7144 6326
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7576 5642 7604 6598
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8312 5370 8340 5578
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 6780 4924 7088 4933
rect 6780 4922 6786 4924
rect 6842 4922 6866 4924
rect 6922 4922 6946 4924
rect 7002 4922 7026 4924
rect 7082 4922 7088 4924
rect 6842 4870 6844 4922
rect 7024 4870 7026 4922
rect 6780 4868 6786 4870
rect 6842 4868 6866 4870
rect 6922 4868 6946 4870
rect 7002 4868 7026 4870
rect 7082 4868 7088 4870
rect 6780 4859 7088 4868
rect 7392 4826 7420 4966
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6656 3738 6684 4082
rect 6780 3836 7088 3845
rect 6780 3834 6786 3836
rect 6842 3834 6866 3836
rect 6922 3834 6946 3836
rect 7002 3834 7026 3836
rect 7082 3834 7088 3836
rect 6842 3782 6844 3834
rect 7024 3782 7026 3834
rect 6780 3780 6786 3782
rect 6842 3780 6866 3782
rect 6922 3780 6946 3782
rect 7002 3780 7026 3782
rect 7082 3780 7088 3782
rect 6780 3771 7088 3780
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 7300 3534 7328 4422
rect 7760 4214 7788 4422
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 3194 7512 3334
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 8312 3058 8340 3402
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 6472 2746 6592 2774
rect 6780 2748 7088 2757
rect 6780 2746 6786 2748
rect 6842 2746 6866 2748
rect 6922 2746 6946 2748
rect 7002 2746 7026 2748
rect 7082 2746 7088 2748
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6472 2446 6500 2746
rect 6842 2694 6844 2746
rect 7024 2694 7026 2746
rect 6780 2692 6786 2694
rect 6842 2692 6866 2694
rect 6922 2692 6946 2694
rect 7002 2692 7026 2694
rect 7082 2692 7088 2694
rect 6780 2683 7088 2692
rect 7116 2650 7144 2994
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7944 2650 7972 2790
rect 8404 2650 8432 10406
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8496 9178 8524 9522
rect 8588 9518 8616 10542
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 8723 9820 9031 9829
rect 8723 9818 8729 9820
rect 8785 9818 8809 9820
rect 8865 9818 8889 9820
rect 8945 9818 8969 9820
rect 9025 9818 9031 9820
rect 8785 9766 8787 9818
rect 8967 9766 8969 9818
rect 8723 9764 8729 9766
rect 8785 9764 8809 9766
rect 8865 9764 8889 9766
rect 8945 9764 8969 9766
rect 9025 9764 9031 9766
rect 8723 9755 9031 9764
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8634 8524 8978
rect 8864 8974 8892 9522
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8634 8616 8774
rect 8723 8732 9031 8741
rect 8723 8730 8729 8732
rect 8785 8730 8809 8732
rect 8865 8730 8889 8732
rect 8945 8730 8969 8732
rect 9025 8730 9031 8732
rect 8785 8678 8787 8730
rect 8967 8678 8969 8730
rect 8723 8676 8729 8678
rect 8785 8676 8809 8678
rect 8865 8676 8889 8678
rect 8945 8676 8969 8678
rect 9025 8676 9031 8678
rect 8723 8667 9031 8676
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9140 8378 9168 10134
rect 9232 8974 9260 11222
rect 9324 9994 9352 11750
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9416 11354 9444 11698
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 10810 9444 11018
rect 9508 10810 9536 12406
rect 9600 11558 9628 14418
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9968 14074 9996 14350
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9956 13184 10008 13190
rect 9692 13144 9956 13172
rect 9692 12434 9720 13144
rect 9956 13126 10008 13132
rect 9862 12744 9918 12753
rect 9862 12679 9918 12688
rect 9692 12406 9812 12434
rect 9784 12238 9812 12406
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11098 9628 11494
rect 9784 11150 9812 11562
rect 9876 11150 9904 12679
rect 10060 12646 10088 15302
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 9772 11144 9824 11150
rect 9600 11070 9720 11098
rect 9772 11086 9824 11092
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9692 10962 9720 11070
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9692 10934 9904 10962
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9508 10690 9536 10746
rect 9416 10662 9536 10690
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9416 10266 9444 10662
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9324 9178 9352 9318
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9232 8498 9260 8910
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 8022 8524 8230
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8496 7206 8524 7958
rect 9048 7886 9076 8366
rect 9140 8350 9260 8378
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8496 2990 8524 7142
rect 8588 3466 8616 7686
rect 8723 7644 9031 7653
rect 8723 7642 8729 7644
rect 8785 7642 8809 7644
rect 8865 7642 8889 7644
rect 8945 7642 8969 7644
rect 9025 7642 9031 7644
rect 8785 7590 8787 7642
rect 8967 7590 8969 7642
rect 8723 7588 8729 7590
rect 8785 7588 8809 7590
rect 8865 7588 8889 7590
rect 8945 7588 8969 7590
rect 9025 7588 9031 7590
rect 8723 7579 9031 7588
rect 8723 6556 9031 6565
rect 8723 6554 8729 6556
rect 8785 6554 8809 6556
rect 8865 6554 8889 6556
rect 8945 6554 8969 6556
rect 9025 6554 9031 6556
rect 8785 6502 8787 6554
rect 8967 6502 8969 6554
rect 8723 6500 8729 6502
rect 8785 6500 8809 6502
rect 8865 6500 8889 6502
rect 8945 6500 8969 6502
rect 9025 6500 9031 6502
rect 8723 6491 9031 6500
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5914 8708 6054
rect 8864 5914 8892 6258
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8723 5468 9031 5477
rect 8723 5466 8729 5468
rect 8785 5466 8809 5468
rect 8865 5466 8889 5468
rect 8945 5466 8969 5468
rect 9025 5466 9031 5468
rect 8785 5414 8787 5466
rect 8967 5414 8969 5466
rect 8723 5412 8729 5414
rect 8785 5412 8809 5414
rect 8865 5412 8889 5414
rect 8945 5412 8969 5414
rect 9025 5412 9031 5414
rect 8723 5403 9031 5412
rect 9232 4622 9260 8350
rect 9324 7818 9352 9114
rect 9416 8616 9444 9862
rect 9508 9518 9536 10542
rect 9692 10266 9720 10678
rect 9784 10606 9812 10746
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9784 10470 9812 10542
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9600 9450 9628 9862
rect 9692 9722 9720 10202
rect 9784 9994 9812 10406
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 9178 9536 9318
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9692 9110 9720 9658
rect 9876 9178 9904 10934
rect 9968 10266 9996 11018
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9416 8588 9536 8616
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 8090 9444 8434
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 5914 9352 6598
rect 9508 6390 9536 8588
rect 9692 8498 9720 9046
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9692 7886 9720 8298
rect 9968 8090 9996 10066
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9968 7290 9996 7754
rect 9876 7262 9996 7290
rect 9876 7206 9904 7262
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6798 9904 7142
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9508 5778 9536 6326
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5370 9628 5510
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 8723 4380 9031 4389
rect 8723 4378 8729 4380
rect 8785 4378 8809 4380
rect 8865 4378 8889 4380
rect 8945 4378 8969 4380
rect 9025 4378 9031 4380
rect 8785 4326 8787 4378
rect 8967 4326 8969 4378
rect 8723 4324 8729 4326
rect 8785 4324 8809 4326
rect 8865 4324 8889 4326
rect 8945 4324 8969 4326
rect 9025 4324 9031 4326
rect 8723 4315 9031 4324
rect 9508 4060 9536 5238
rect 9600 4486 9628 5306
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9784 4826 9812 5170
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9588 4072 9640 4078
rect 9508 4032 9588 4060
rect 9588 4014 9640 4020
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8723 3292 9031 3301
rect 8723 3290 8729 3292
rect 8785 3290 8809 3292
rect 8865 3290 8889 3292
rect 8945 3290 8969 3292
rect 9025 3290 9031 3292
rect 8785 3238 8787 3290
rect 8967 3238 8969 3290
rect 8723 3236 8729 3238
rect 8785 3236 8809 3238
rect 8865 3236 8889 3238
rect 8945 3236 8969 3238
rect 9025 3236 9031 3238
rect 8723 3227 9031 3236
rect 9600 3126 9628 4014
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 10060 2446 10088 12582
rect 10152 10674 10180 17002
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 10667 16892 10975 16901
rect 10667 16890 10673 16892
rect 10729 16890 10753 16892
rect 10809 16890 10833 16892
rect 10889 16890 10913 16892
rect 10969 16890 10975 16892
rect 10729 16838 10731 16890
rect 10911 16838 10913 16890
rect 10667 16836 10673 16838
rect 10729 16836 10753 16838
rect 10809 16836 10833 16838
rect 10889 16836 10913 16838
rect 10969 16836 10975 16838
rect 10667 16827 10975 16836
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10244 12986 10272 15574
rect 10428 15434 10456 16050
rect 10667 15804 10975 15813
rect 10667 15802 10673 15804
rect 10729 15802 10753 15804
rect 10809 15802 10833 15804
rect 10889 15802 10913 15804
rect 10969 15802 10975 15804
rect 10729 15750 10731 15802
rect 10911 15750 10913 15802
rect 10667 15748 10673 15750
rect 10729 15748 10753 15750
rect 10809 15748 10833 15750
rect 10889 15748 10913 15750
rect 10969 15748 10975 15750
rect 10667 15739 10975 15748
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10428 14550 10456 15370
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10520 14618 10548 15030
rect 10667 14716 10975 14725
rect 10667 14714 10673 14716
rect 10729 14714 10753 14716
rect 10809 14714 10833 14716
rect 10889 14714 10913 14716
rect 10969 14714 10975 14716
rect 10729 14662 10731 14714
rect 10911 14662 10913 14714
rect 10667 14660 10673 14662
rect 10729 14660 10753 14662
rect 10809 14660 10833 14662
rect 10889 14660 10913 14662
rect 10969 14660 10975 14662
rect 10667 14651 10975 14660
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10336 13530 10364 13874
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10232 12980 10284 12986
rect 10284 12940 10364 12968
rect 10232 12922 10284 12928
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10244 12102 10272 12786
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10244 11626 10272 12038
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10152 10470 10180 10610
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 9042 10180 10406
rect 10336 10130 10364 12940
rect 10428 12918 10456 14486
rect 11072 14482 11100 16594
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11348 14958 11376 16050
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11532 15094 11560 15982
rect 11900 15638 11928 16934
rect 14554 16892 14862 16901
rect 14554 16890 14560 16892
rect 14616 16890 14640 16892
rect 14696 16890 14720 16892
rect 14776 16890 14800 16892
rect 14856 16890 14862 16892
rect 14616 16838 14618 16890
rect 14798 16838 14800 16890
rect 14554 16836 14560 16838
rect 14616 16836 14640 16838
rect 14696 16836 14720 16838
rect 14776 16836 14800 16838
rect 14856 16836 14862 16838
rect 14554 16827 14862 16836
rect 12610 16348 12918 16357
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12268 15706 12296 16118
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 13096 15094 13124 15302
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10520 11234 10548 14214
rect 11072 14090 11100 14418
rect 11072 14062 11192 14090
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10667 13628 10975 13637
rect 10667 13626 10673 13628
rect 10729 13626 10753 13628
rect 10809 13626 10833 13628
rect 10889 13626 10913 13628
rect 10969 13626 10975 13628
rect 10729 13574 10731 13626
rect 10911 13574 10913 13626
rect 10667 13572 10673 13574
rect 10729 13572 10753 13574
rect 10809 13572 10833 13574
rect 10889 13572 10913 13574
rect 10969 13572 10975 13574
rect 10667 13563 10975 13572
rect 11072 13530 11100 13874
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 11072 12918 11100 13466
rect 11164 13190 11192 14062
rect 11256 13802 11284 14894
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11440 13326 11468 13942
rect 11532 13938 11560 14282
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11348 12986 11376 13194
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10667 12540 10975 12549
rect 10667 12538 10673 12540
rect 10729 12538 10753 12540
rect 10809 12538 10833 12540
rect 10889 12538 10913 12540
rect 10969 12538 10975 12540
rect 10729 12486 10731 12538
rect 10911 12486 10913 12538
rect 10667 12484 10673 12486
rect 10729 12484 10753 12486
rect 10809 12484 10833 12486
rect 10889 12484 10913 12486
rect 10969 12484 10975 12486
rect 10667 12475 10975 12484
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 10667 11452 10975 11461
rect 10667 11450 10673 11452
rect 10729 11450 10753 11452
rect 10809 11450 10833 11452
rect 10889 11450 10913 11452
rect 10969 11450 10975 11452
rect 10729 11398 10731 11450
rect 10911 11398 10913 11450
rect 10667 11396 10673 11398
rect 10729 11396 10753 11398
rect 10809 11396 10833 11398
rect 10889 11396 10913 11398
rect 10969 11396 10975 11398
rect 10667 11387 10975 11396
rect 10520 11206 10640 11234
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10152 8498 10180 8978
rect 10244 8974 10272 9318
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10336 8430 10364 9454
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10428 8362 10456 9522
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7546 10272 7686
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10520 6798 10548 11086
rect 10612 10742 10640 11206
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10667 10364 10975 10373
rect 10667 10362 10673 10364
rect 10729 10362 10753 10364
rect 10809 10362 10833 10364
rect 10889 10362 10913 10364
rect 10969 10362 10975 10364
rect 10729 10310 10731 10362
rect 10911 10310 10913 10362
rect 10667 10308 10673 10310
rect 10729 10308 10753 10310
rect 10809 10308 10833 10310
rect 10889 10308 10913 10310
rect 10969 10308 10975 10310
rect 10667 10299 10975 10308
rect 10667 9276 10975 9285
rect 10667 9274 10673 9276
rect 10729 9274 10753 9276
rect 10809 9274 10833 9276
rect 10889 9274 10913 9276
rect 10969 9274 10975 9276
rect 10729 9222 10731 9274
rect 10911 9222 10913 9274
rect 10667 9220 10673 9222
rect 10729 9220 10753 9222
rect 10809 9220 10833 9222
rect 10889 9220 10913 9222
rect 10969 9220 10975 9222
rect 10667 9211 10975 9220
rect 11072 9042 11100 10610
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11164 9586 11192 10202
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11256 9178 11284 9998
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11072 8498 11100 8978
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10667 8188 10975 8197
rect 10667 8186 10673 8188
rect 10729 8186 10753 8188
rect 10809 8186 10833 8188
rect 10889 8186 10913 8188
rect 10969 8186 10975 8188
rect 10729 8134 10731 8186
rect 10911 8134 10913 8186
rect 10667 8132 10673 8134
rect 10729 8132 10753 8134
rect 10809 8132 10833 8134
rect 10889 8132 10913 8134
rect 10969 8132 10975 8134
rect 10667 8123 10975 8132
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10980 7886 11008 8026
rect 11072 8022 11100 8298
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10667 7100 10975 7109
rect 10667 7098 10673 7100
rect 10729 7098 10753 7100
rect 10809 7098 10833 7100
rect 10889 7098 10913 7100
rect 10969 7098 10975 7100
rect 10729 7046 10731 7098
rect 10911 7046 10913 7098
rect 10667 7044 10673 7046
rect 10729 7044 10753 7046
rect 10809 7044 10833 7046
rect 10889 7044 10913 7046
rect 10969 7044 10975 7046
rect 10667 7035 10975 7044
rect 11072 7002 11100 7346
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 11164 6662 11192 7686
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 11256 6798 11284 6870
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11348 6322 11376 11698
rect 11440 7290 11468 13262
rect 11532 12434 11560 13874
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11808 12434 11836 12854
rect 11900 12850 11928 13194
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11532 12406 11652 12434
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11532 8634 11560 8842
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11440 7262 11560 7290
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 6730 11468 7142
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 10667 6012 10975 6021
rect 10667 6010 10673 6012
rect 10729 6010 10753 6012
rect 10809 6010 10833 6012
rect 10889 6010 10913 6012
rect 10969 6010 10975 6012
rect 10729 5958 10731 6010
rect 10911 5958 10913 6010
rect 10667 5956 10673 5958
rect 10729 5956 10753 5958
rect 10809 5956 10833 5958
rect 10889 5956 10913 5958
rect 10969 5956 10975 5958
rect 10667 5947 10975 5956
rect 11440 5778 11468 6666
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10428 5370 10456 5578
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 11532 5114 11560 7262
rect 11624 5234 11652 12406
rect 11716 12406 11836 12434
rect 11716 11830 11744 12406
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11716 11150 11744 11766
rect 11900 11762 11928 12786
rect 11992 12442 12020 14894
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12084 12918 12112 13806
rect 12176 13258 12204 13874
rect 12268 13870 12296 15030
rect 13188 14618 13216 15982
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 15706 13400 15846
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13740 14958 13768 15914
rect 14554 15804 14862 15813
rect 14554 15802 14560 15804
rect 14616 15802 14640 15804
rect 14696 15802 14720 15804
rect 14776 15802 14800 15804
rect 14856 15802 14862 15804
rect 14616 15750 14618 15802
rect 14798 15750 14800 15802
rect 14554 15748 14560 15750
rect 14616 15748 14640 15750
rect 14696 15748 14720 15750
rect 14776 15748 14800 15750
rect 14856 15748 14862 15750
rect 14554 15739 14862 15748
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14200 15094 14228 15302
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12360 14074 12388 14282
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 13188 14074 13216 14554
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 13004 13530 13032 13874
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12176 12782 12204 13194
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12986 12480 13126
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11992 11830 12020 12378
rect 12544 12238 12572 12582
rect 13372 12442 13400 12854
rect 13648 12850 13676 14758
rect 13740 14482 13768 14894
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13740 12918 13768 14418
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14108 14074 14136 14214
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14292 13734 14320 14214
rect 14384 14074 14412 15438
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14476 14414 14504 14758
rect 14554 14716 14862 14725
rect 14554 14714 14560 14716
rect 14616 14714 14640 14716
rect 14696 14714 14720 14716
rect 14776 14714 14800 14716
rect 14856 14714 14862 14716
rect 14616 14662 14618 14714
rect 14798 14662 14800 14714
rect 14554 14660 14560 14662
rect 14616 14660 14640 14662
rect 14696 14660 14720 14662
rect 14776 14660 14800 14662
rect 14856 14660 14862 14662
rect 14554 14651 14862 14660
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 13832 13394 13860 13670
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13832 12918 13860 13330
rect 14292 13258 14320 13670
rect 14384 13394 14412 13738
rect 14554 13628 14862 13637
rect 14554 13626 14560 13628
rect 14616 13626 14640 13628
rect 14696 13626 14720 13628
rect 14776 13626 14800 13628
rect 14856 13626 14862 13628
rect 14616 13574 14618 13626
rect 14798 13574 14800 13626
rect 14554 13572 14560 13574
rect 14616 13572 14640 13574
rect 14696 13572 14720 13574
rect 14776 13572 14800 13574
rect 14856 13572 14862 13574
rect 14554 13563 14862 13572
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 15396 13258 15424 13942
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13832 12238 13860 12582
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12084 11898 12112 12106
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 12268 11762 12296 12174
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 11900 11218 11928 11698
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11716 10810 11744 11086
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11900 10266 11928 11154
rect 12268 11150 12296 11698
rect 12256 11144 12308 11150
rect 12308 11092 12480 11098
rect 12256 11086 12480 11092
rect 12268 11070 12480 11086
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 12084 10062 12112 10746
rect 12452 10130 12480 11070
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12610 10843 12918 10852
rect 13924 10674 13952 12718
rect 14554 12540 14862 12549
rect 14554 12538 14560 12540
rect 14616 12538 14640 12540
rect 14696 12538 14720 12540
rect 14776 12538 14800 12540
rect 14856 12538 14862 12540
rect 14616 12486 14618 12538
rect 14798 12486 14800 12538
rect 14554 12484 14560 12486
rect 14616 12484 14640 12486
rect 14696 12484 14720 12486
rect 14776 12484 14800 12486
rect 14856 12484 14862 12486
rect 14554 12475 14862 12484
rect 15764 12170 15792 16934
rect 16497 16348 16805 16357
rect 16497 16346 16503 16348
rect 16559 16346 16583 16348
rect 16639 16346 16663 16348
rect 16719 16346 16743 16348
rect 16799 16346 16805 16348
rect 16559 16294 16561 16346
rect 16741 16294 16743 16346
rect 16497 16292 16503 16294
rect 16559 16292 16583 16294
rect 16639 16292 16663 16294
rect 16719 16292 16743 16294
rect 16799 16292 16805 16294
rect 16497 16283 16805 16292
rect 16497 15260 16805 15269
rect 16497 15258 16503 15260
rect 16559 15258 16583 15260
rect 16639 15258 16663 15260
rect 16719 15258 16743 15260
rect 16799 15258 16805 15260
rect 16559 15206 16561 15258
rect 16741 15206 16743 15258
rect 16497 15204 16503 15206
rect 16559 15204 16583 15206
rect 16639 15204 16663 15206
rect 16719 15204 16743 15206
rect 16799 15204 16805 15206
rect 16497 15195 16805 15204
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16224 14074 16252 14214
rect 16497 14172 16805 14181
rect 16497 14170 16503 14172
rect 16559 14170 16583 14172
rect 16639 14170 16663 14172
rect 16719 14170 16743 14172
rect 16799 14170 16805 14172
rect 16559 14118 16561 14170
rect 16741 14118 16743 14170
rect 16497 14116 16503 14118
rect 16559 14116 16583 14118
rect 16639 14116 16663 14118
rect 16719 14116 16743 14118
rect 16799 14116 16805 14118
rect 16497 14107 16805 14116
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16592 13705 16620 13806
rect 16578 13696 16634 13705
rect 16578 13631 16634 13640
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12986 15884 13126
rect 16497 13084 16805 13093
rect 16497 13082 16503 13084
rect 16559 13082 16583 13084
rect 16639 13082 16663 13084
rect 16719 13082 16743 13084
rect 16799 13082 16805 13084
rect 16559 13030 16561 13082
rect 16741 13030 16743 13082
rect 16497 13028 16503 13030
rect 16559 13028 16583 13030
rect 16639 13028 16663 13030
rect 16719 13028 16743 13030
rect 16799 13028 16805 13030
rect 16497 13019 16805 13028
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15752 12164 15804 12170
rect 15752 12106 15804 12112
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14108 11898 14136 12038
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 14554 11452 14862 11461
rect 14554 11450 14560 11452
rect 14616 11450 14640 11452
rect 14696 11450 14720 11452
rect 14776 11450 14800 11452
rect 14856 11450 14862 11452
rect 14616 11398 14618 11450
rect 14798 11398 14800 11450
rect 14554 11396 14560 11398
rect 14616 11396 14640 11398
rect 14696 11396 14720 11398
rect 14776 11396 14800 11398
rect 14856 11396 14862 11398
rect 14554 11387 14862 11396
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14292 10810 14320 11290
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 13740 10062 13768 10406
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 12084 9722 12112 9998
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 13924 9722 13952 10202
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 11888 9376 11940 9382
rect 11940 9324 12020 9330
rect 11888 9318 12020 9324
rect 11900 9302 12020 9318
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11808 7970 11836 8298
rect 11900 8090 11928 8774
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11808 7942 11928 7970
rect 11900 7886 11928 7942
rect 11992 7886 12020 9302
rect 12912 9178 12940 9386
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8634 12572 8774
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11900 6934 11928 7822
rect 11992 7206 12020 7822
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 7546 12112 7686
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11992 6866 12020 7142
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6322 11836 6598
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11808 5234 11836 6258
rect 12084 5846 12112 7346
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12176 6322 12204 6870
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11992 5370 12020 5510
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12084 5302 12112 5782
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11532 5086 11744 5114
rect 10667 4924 10975 4933
rect 10667 4922 10673 4924
rect 10729 4922 10753 4924
rect 10809 4922 10833 4924
rect 10889 4922 10913 4924
rect 10969 4922 10975 4924
rect 10729 4870 10731 4922
rect 10911 4870 10913 4922
rect 10667 4868 10673 4870
rect 10729 4868 10753 4870
rect 10809 4868 10833 4870
rect 10889 4868 10913 4870
rect 10969 4868 10975 4870
rect 10667 4859 10975 4868
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10152 4214 10180 4422
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10336 3738 10364 4558
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10667 3836 10975 3845
rect 10667 3834 10673 3836
rect 10729 3834 10753 3836
rect 10809 3834 10833 3836
rect 10889 3834 10913 3836
rect 10969 3834 10975 3836
rect 10729 3782 10731 3834
rect 10911 3782 10913 3834
rect 10667 3780 10673 3782
rect 10729 3780 10753 3782
rect 10809 3780 10833 3782
rect 10889 3780 10913 3782
rect 10969 3780 10975 3782
rect 10667 3771 10975 3780
rect 11072 3738 11100 3946
rect 11532 3738 11560 4082
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6460 2440 6512 2446
rect 7840 2440 7892 2446
rect 6460 2382 6512 2388
rect 7760 2400 7840 2428
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 4836 2204 5144 2213
rect 4836 2202 4842 2204
rect 4898 2202 4922 2204
rect 4978 2202 5002 2204
rect 5058 2202 5082 2204
rect 5138 2202 5144 2204
rect 4898 2150 4900 2202
rect 5080 2150 5082 2202
rect 4836 2148 4842 2150
rect 4898 2148 4922 2150
rect 4978 2148 5002 2150
rect 5058 2148 5082 2150
rect 5138 2148 5144 2150
rect 4836 2139 5144 2148
rect 3896 1142 4108 1170
rect 3896 800 3924 1142
rect 7760 800 7788 2400
rect 7840 2382 7892 2388
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10428 2378 10456 2790
rect 10520 2650 10548 2994
rect 10796 2854 10824 3334
rect 11716 3194 11744 5086
rect 11808 4622 11836 5170
rect 12084 4706 12112 5238
rect 12176 5234 12204 6258
rect 12268 5914 12296 6258
rect 12360 6254 12388 6802
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 11900 4678 12112 4706
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10667 2748 10975 2757
rect 10667 2746 10673 2748
rect 10729 2746 10753 2748
rect 10809 2746 10833 2748
rect 10889 2746 10913 2748
rect 10969 2746 10975 2748
rect 10729 2694 10731 2746
rect 10911 2694 10913 2746
rect 10667 2692 10673 2694
rect 10729 2692 10753 2694
rect 10809 2692 10833 2694
rect 10889 2692 10913 2694
rect 10969 2692 10975 2694
rect 10667 2683 10975 2692
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 11716 2582 11744 3130
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 10416 2372 10468 2378
rect 10416 2314 10468 2320
rect 11808 2310 11836 4558
rect 11900 3602 11928 4678
rect 12176 4622 12204 5170
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11900 3058 11928 3538
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11900 2514 12020 2530
rect 11900 2508 12032 2514
rect 11900 2502 11980 2508
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 8723 2204 9031 2213
rect 8723 2202 8729 2204
rect 8785 2202 8809 2204
rect 8865 2202 8889 2204
rect 8945 2202 8969 2204
rect 9025 2202 9031 2204
rect 8785 2150 8787 2202
rect 8967 2150 8969 2202
rect 8723 2148 8729 2150
rect 8785 2148 8809 2150
rect 8865 2148 8889 2150
rect 8945 2148 8969 2150
rect 9025 2148 9031 2150
rect 8723 2139 9031 2148
rect 11624 870 11744 898
rect 11624 800 11652 870
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 11716 762 11744 870
rect 11900 762 11928 2502
rect 11980 2450 12032 2456
rect 12176 2446 12204 4558
rect 12268 4146 12296 5850
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12360 4146 12388 5510
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12268 3602 12296 3878
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12268 2650 12296 2994
rect 12452 2650 12480 8366
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12544 7954 12572 8230
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 13740 7546 13768 7754
rect 13832 7546 13860 7822
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 13648 5710 13676 7346
rect 13924 6866 13952 8910
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7546 14136 7686
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 7002 14044 7142
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14292 6730 14320 10610
rect 14554 10364 14862 10373
rect 14554 10362 14560 10364
rect 14616 10362 14640 10364
rect 14696 10362 14720 10364
rect 14776 10362 14800 10364
rect 14856 10362 14862 10364
rect 14616 10310 14618 10362
rect 14798 10310 14800 10362
rect 14554 10308 14560 10310
rect 14616 10308 14640 10310
rect 14696 10308 14720 10310
rect 14776 10308 14800 10310
rect 14856 10308 14862 10310
rect 14554 10299 14862 10308
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14568 9722 14596 9862
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14936 9518 14964 11154
rect 15028 10810 15056 11766
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 11354 15516 11494
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15764 11286 15792 12106
rect 16497 11996 16805 12005
rect 16497 11994 16503 11996
rect 16559 11994 16583 11996
rect 16639 11994 16663 11996
rect 16719 11994 16743 11996
rect 16799 11994 16805 11996
rect 16559 11942 16561 11994
rect 16741 11942 16743 11994
rect 16497 11940 16503 11942
rect 16559 11940 16583 11942
rect 16639 11940 16663 11942
rect 16719 11940 16743 11942
rect 16799 11940 16805 11942
rect 16497 11931 16805 11940
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15856 11354 15884 11630
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15212 10810 15240 11222
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 15028 9654 15056 10610
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15120 10130 15148 10406
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15396 9722 15424 9930
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 15028 9466 15056 9590
rect 14554 9276 14862 9285
rect 14554 9274 14560 9276
rect 14616 9274 14640 9276
rect 14696 9274 14720 9276
rect 14776 9274 14800 9276
rect 14856 9274 14862 9276
rect 14616 9222 14618 9274
rect 14798 9222 14800 9274
rect 14554 9220 14560 9222
rect 14616 9220 14640 9222
rect 14696 9220 14720 9222
rect 14776 9220 14800 9222
rect 14856 9220 14862 9222
rect 14554 9211 14862 9220
rect 14936 9178 14964 9454
rect 15028 9438 15148 9466
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14554 8188 14862 8197
rect 14554 8186 14560 8188
rect 14616 8186 14640 8188
rect 14696 8186 14720 8188
rect 14776 8186 14800 8188
rect 14856 8186 14862 8188
rect 14616 8134 14618 8186
rect 14798 8134 14800 8186
rect 14554 8132 14560 8134
rect 14616 8132 14640 8134
rect 14696 8132 14720 8134
rect 14776 8132 14800 8134
rect 14856 8132 14862 8134
rect 14554 8123 14862 8132
rect 14936 7954 14964 9114
rect 15028 9042 15056 9318
rect 15120 9042 15148 9438
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 14554 7100 14862 7109
rect 14554 7098 14560 7100
rect 14616 7098 14640 7100
rect 14696 7098 14720 7100
rect 14776 7098 14800 7100
rect 14856 7098 14862 7100
rect 14616 7046 14618 7098
rect 14798 7046 14800 7098
rect 14554 7044 14560 7046
rect 14616 7044 14640 7046
rect 14696 7044 14720 7046
rect 14776 7044 14800 7046
rect 14856 7044 14862 7046
rect 14554 7035 14862 7044
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14292 6202 14320 6666
rect 14936 6254 14964 7890
rect 15120 7478 15148 8978
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 6730 15424 7142
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 14200 6174 14320 6202
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 12636 5556 12664 5646
rect 12544 5528 12664 5556
rect 12544 3738 12572 5528
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4826 13676 4966
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 13176 4072 13228 4078
rect 13832 4026 13860 4694
rect 13924 4214 13952 5170
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 13176 4014 13228 4020
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 13188 3194 13216 4014
rect 13740 4010 13860 4026
rect 13728 4004 13860 4010
rect 13780 3998 13860 4004
rect 13728 3946 13780 3952
rect 13924 3738 13952 4150
rect 14016 4078 14044 4422
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 14200 3670 14228 6174
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14292 5914 14320 6054
rect 14554 6012 14862 6021
rect 14554 6010 14560 6012
rect 14616 6010 14640 6012
rect 14696 6010 14720 6012
rect 14776 6010 14800 6012
rect 14856 6010 14862 6012
rect 14616 5958 14618 6010
rect 14798 5958 14800 6010
rect 14554 5956 14560 5958
rect 14616 5956 14640 5958
rect 14696 5956 14720 5958
rect 14776 5956 14800 5958
rect 14856 5956 14862 5958
rect 14554 5947 14862 5956
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14384 5302 14412 5510
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14554 4924 14862 4933
rect 14554 4922 14560 4924
rect 14616 4922 14640 4924
rect 14696 4922 14720 4924
rect 14776 4922 14800 4924
rect 14856 4922 14862 4924
rect 14616 4870 14618 4922
rect 14798 4870 14800 4922
rect 14554 4868 14560 4870
rect 14616 4868 14640 4870
rect 14696 4868 14720 4870
rect 14776 4868 14800 4870
rect 14856 4868 14862 4870
rect 14554 4859 14862 4868
rect 14936 4690 14964 6190
rect 15764 5234 15792 7346
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15856 6458 15884 6598
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 16132 5914 16160 11018
rect 16497 10908 16805 10917
rect 16497 10906 16503 10908
rect 16559 10906 16583 10908
rect 16639 10906 16663 10908
rect 16719 10906 16743 10908
rect 16799 10906 16805 10908
rect 16559 10854 16561 10906
rect 16741 10854 16743 10906
rect 16497 10852 16503 10854
rect 16559 10852 16583 10854
rect 16639 10852 16663 10854
rect 16719 10852 16743 10854
rect 16799 10852 16805 10854
rect 16497 10843 16805 10852
rect 16497 9820 16805 9829
rect 16497 9818 16503 9820
rect 16559 9818 16583 9820
rect 16639 9818 16663 9820
rect 16719 9818 16743 9820
rect 16799 9818 16805 9820
rect 16559 9766 16561 9818
rect 16741 9766 16743 9818
rect 16497 9764 16503 9766
rect 16559 9764 16583 9766
rect 16639 9764 16663 9766
rect 16719 9764 16743 9766
rect 16799 9764 16805 9766
rect 16497 9755 16805 9764
rect 16302 9616 16358 9625
rect 16302 9551 16304 9560
rect 16356 9551 16358 9560
rect 16304 9522 16356 9528
rect 16497 8732 16805 8741
rect 16497 8730 16503 8732
rect 16559 8730 16583 8732
rect 16639 8730 16663 8732
rect 16719 8730 16743 8732
rect 16799 8730 16805 8732
rect 16559 8678 16561 8730
rect 16741 8678 16743 8730
rect 16497 8676 16503 8678
rect 16559 8676 16583 8678
rect 16639 8676 16663 8678
rect 16719 8676 16743 8678
rect 16799 8676 16805 8678
rect 16497 8667 16805 8676
rect 16497 7644 16805 7653
rect 16497 7642 16503 7644
rect 16559 7642 16583 7644
rect 16639 7642 16663 7644
rect 16719 7642 16743 7644
rect 16799 7642 16805 7644
rect 16559 7590 16561 7642
rect 16741 7590 16743 7642
rect 16497 7588 16503 7590
rect 16559 7588 16583 7590
rect 16639 7588 16663 7590
rect 16719 7588 16743 7590
rect 16799 7588 16805 7590
rect 16497 7579 16805 7588
rect 16497 6556 16805 6565
rect 16497 6554 16503 6556
rect 16559 6554 16583 6556
rect 16639 6554 16663 6556
rect 16719 6554 16743 6556
rect 16799 6554 16805 6556
rect 16559 6502 16561 6554
rect 16741 6502 16743 6554
rect 16497 6500 16503 6502
rect 16559 6500 16583 6502
rect 16639 6500 16663 6502
rect 16719 6500 16743 6502
rect 16799 6500 16805 6502
rect 16497 6491 16805 6500
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 16960 5545 16988 5578
rect 16946 5536 17002 5545
rect 16497 5468 16805 5477
rect 16946 5471 17002 5480
rect 16497 5466 16503 5468
rect 16559 5466 16583 5468
rect 16639 5466 16663 5468
rect 16719 5466 16743 5468
rect 16799 5466 16805 5468
rect 16559 5414 16561 5466
rect 16741 5414 16743 5466
rect 16497 5412 16503 5414
rect 16559 5412 16583 5414
rect 16639 5412 16663 5414
rect 16719 5412 16743 5414
rect 16799 5412 16805 5414
rect 16497 5403 16805 5412
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 15764 4078 15792 5170
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 4826 15976 4966
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 16497 4380 16805 4389
rect 16497 4378 16503 4380
rect 16559 4378 16583 4380
rect 16639 4378 16663 4380
rect 16719 4378 16743 4380
rect 16799 4378 16805 4380
rect 16559 4326 16561 4378
rect 16741 4326 16743 4378
rect 16497 4324 16503 4326
rect 16559 4324 16583 4326
rect 16639 4324 16663 4326
rect 16719 4324 16743 4326
rect 16799 4324 16805 4326
rect 16497 4315 16805 4324
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 14554 3836 14862 3845
rect 14554 3834 14560 3836
rect 14616 3834 14640 3836
rect 14696 3834 14720 3836
rect 14776 3834 14800 3836
rect 14856 3834 14862 3836
rect 14616 3782 14618 3834
rect 14798 3782 14800 3834
rect 14554 3780 14560 3782
rect 14616 3780 14640 3782
rect 14696 3780 14720 3782
rect 14776 3780 14800 3782
rect 14856 3780 14862 3782
rect 14554 3771 14862 3780
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13188 2774 13216 3130
rect 13188 2746 13400 2774
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 13372 2378 13400 2746
rect 14554 2748 14862 2757
rect 14554 2746 14560 2748
rect 14616 2746 14640 2748
rect 14696 2746 14720 2748
rect 14776 2746 14800 2748
rect 14856 2746 14862 2748
rect 14616 2694 14618 2746
rect 14798 2694 14800 2746
rect 14554 2692 14560 2694
rect 14616 2692 14640 2694
rect 14696 2692 14720 2694
rect 14776 2692 14800 2694
rect 14856 2692 14862 2694
rect 14554 2683 14862 2692
rect 16132 2650 16160 3402
rect 16497 3292 16805 3301
rect 16497 3290 16503 3292
rect 16559 3290 16583 3292
rect 16639 3290 16663 3292
rect 16719 3290 16743 3292
rect 16799 3290 16805 3292
rect 16559 3238 16561 3290
rect 16741 3238 16743 3290
rect 16497 3236 16503 3238
rect 16559 3236 16583 3238
rect 16639 3236 16663 3238
rect 16719 3236 16743 3238
rect 16799 3236 16805 3238
rect 16497 3227 16805 3236
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 15672 1170 15700 2314
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16408 1442 16436 2246
rect 16497 2204 16805 2213
rect 16497 2202 16503 2204
rect 16559 2202 16583 2204
rect 16639 2202 16663 2204
rect 16719 2202 16743 2204
rect 16799 2202 16805 2204
rect 16559 2150 16561 2202
rect 16741 2150 16743 2202
rect 16497 2148 16503 2150
rect 16559 2148 16583 2150
rect 16639 2148 16663 2150
rect 16719 2148 16743 2150
rect 16799 2148 16805 2150
rect 16497 2139 16805 2148
rect 16486 1456 16542 1465
rect 16408 1414 16486 1442
rect 16486 1391 16542 1400
rect 15488 1142 15700 1170
rect 15488 800 15516 1142
rect 11716 734 11928 762
rect 15474 0 15530 800
<< via2 >>
rect 4842 17434 4898 17436
rect 4922 17434 4978 17436
rect 5002 17434 5058 17436
rect 5082 17434 5138 17436
rect 4842 17382 4888 17434
rect 4888 17382 4898 17434
rect 4922 17382 4952 17434
rect 4952 17382 4964 17434
rect 4964 17382 4978 17434
rect 5002 17382 5016 17434
rect 5016 17382 5028 17434
rect 5028 17382 5058 17434
rect 5082 17382 5092 17434
rect 5092 17382 5138 17434
rect 4842 17380 4898 17382
rect 4922 17380 4978 17382
rect 5002 17380 5058 17382
rect 5082 17380 5138 17382
rect 938 16360 994 16416
rect 2899 16890 2955 16892
rect 2979 16890 3035 16892
rect 3059 16890 3115 16892
rect 3139 16890 3195 16892
rect 2899 16838 2945 16890
rect 2945 16838 2955 16890
rect 2979 16838 3009 16890
rect 3009 16838 3021 16890
rect 3021 16838 3035 16890
rect 3059 16838 3073 16890
rect 3073 16838 3085 16890
rect 3085 16838 3115 16890
rect 3139 16838 3149 16890
rect 3149 16838 3195 16890
rect 2899 16836 2955 16838
rect 2979 16836 3035 16838
rect 3059 16836 3115 16838
rect 3139 16836 3195 16838
rect 1582 12280 1638 12336
rect 2899 15802 2955 15804
rect 2979 15802 3035 15804
rect 3059 15802 3115 15804
rect 3139 15802 3195 15804
rect 2899 15750 2945 15802
rect 2945 15750 2955 15802
rect 2979 15750 3009 15802
rect 3009 15750 3021 15802
rect 3021 15750 3035 15802
rect 3059 15750 3073 15802
rect 3073 15750 3085 15802
rect 3085 15750 3115 15802
rect 3139 15750 3149 15802
rect 3149 15750 3195 15802
rect 2899 15748 2955 15750
rect 2979 15748 3035 15750
rect 3059 15748 3115 15750
rect 3139 15748 3195 15750
rect 2899 14714 2955 14716
rect 2979 14714 3035 14716
rect 3059 14714 3115 14716
rect 3139 14714 3195 14716
rect 2899 14662 2945 14714
rect 2945 14662 2955 14714
rect 2979 14662 3009 14714
rect 3009 14662 3021 14714
rect 3021 14662 3035 14714
rect 3059 14662 3073 14714
rect 3073 14662 3085 14714
rect 3085 14662 3115 14714
rect 3139 14662 3149 14714
rect 3149 14662 3195 14714
rect 2899 14660 2955 14662
rect 2979 14660 3035 14662
rect 3059 14660 3115 14662
rect 3139 14660 3195 14662
rect 2899 13626 2955 13628
rect 2979 13626 3035 13628
rect 3059 13626 3115 13628
rect 3139 13626 3195 13628
rect 2899 13574 2945 13626
rect 2945 13574 2955 13626
rect 2979 13574 3009 13626
rect 3009 13574 3021 13626
rect 3021 13574 3035 13626
rect 3059 13574 3073 13626
rect 3073 13574 3085 13626
rect 3085 13574 3115 13626
rect 3139 13574 3149 13626
rect 3149 13574 3195 13626
rect 2899 13572 2955 13574
rect 2979 13572 3035 13574
rect 3059 13572 3115 13574
rect 3139 13572 3195 13574
rect 8729 17434 8785 17436
rect 8809 17434 8865 17436
rect 8889 17434 8945 17436
rect 8969 17434 9025 17436
rect 8729 17382 8775 17434
rect 8775 17382 8785 17434
rect 8809 17382 8839 17434
rect 8839 17382 8851 17434
rect 8851 17382 8865 17434
rect 8889 17382 8903 17434
rect 8903 17382 8915 17434
rect 8915 17382 8945 17434
rect 8969 17382 8979 17434
rect 8979 17382 9025 17434
rect 8729 17380 8785 17382
rect 8809 17380 8865 17382
rect 8889 17380 8945 17382
rect 8969 17380 9025 17382
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 15934 17720 15990 17776
rect 16503 17434 16559 17436
rect 16583 17434 16639 17436
rect 16663 17434 16719 17436
rect 16743 17434 16799 17436
rect 16503 17382 16549 17434
rect 16549 17382 16559 17434
rect 16583 17382 16613 17434
rect 16613 17382 16625 17434
rect 16625 17382 16639 17434
rect 16663 17382 16677 17434
rect 16677 17382 16689 17434
rect 16689 17382 16719 17434
rect 16743 17382 16753 17434
rect 16753 17382 16799 17434
rect 16503 17380 16559 17382
rect 16583 17380 16639 17382
rect 16663 17380 16719 17382
rect 16743 17380 16799 17382
rect 4842 16346 4898 16348
rect 4922 16346 4978 16348
rect 5002 16346 5058 16348
rect 5082 16346 5138 16348
rect 4842 16294 4888 16346
rect 4888 16294 4898 16346
rect 4922 16294 4952 16346
rect 4952 16294 4964 16346
rect 4964 16294 4978 16346
rect 5002 16294 5016 16346
rect 5016 16294 5028 16346
rect 5028 16294 5058 16346
rect 5082 16294 5092 16346
rect 5092 16294 5138 16346
rect 4842 16292 4898 16294
rect 4922 16292 4978 16294
rect 5002 16292 5058 16294
rect 5082 16292 5138 16294
rect 6786 16890 6842 16892
rect 6866 16890 6922 16892
rect 6946 16890 7002 16892
rect 7026 16890 7082 16892
rect 6786 16838 6832 16890
rect 6832 16838 6842 16890
rect 6866 16838 6896 16890
rect 6896 16838 6908 16890
rect 6908 16838 6922 16890
rect 6946 16838 6960 16890
rect 6960 16838 6972 16890
rect 6972 16838 7002 16890
rect 7026 16838 7036 16890
rect 7036 16838 7082 16890
rect 6786 16836 6842 16838
rect 6866 16836 6922 16838
rect 6946 16836 7002 16838
rect 7026 16836 7082 16838
rect 2899 12538 2955 12540
rect 2979 12538 3035 12540
rect 3059 12538 3115 12540
rect 3139 12538 3195 12540
rect 2899 12486 2945 12538
rect 2945 12486 2955 12538
rect 2979 12486 3009 12538
rect 3009 12486 3021 12538
rect 3021 12486 3035 12538
rect 3059 12486 3073 12538
rect 3073 12486 3085 12538
rect 3085 12486 3115 12538
rect 3139 12486 3149 12538
rect 3149 12486 3195 12538
rect 2899 12484 2955 12486
rect 2979 12484 3035 12486
rect 3059 12484 3115 12486
rect 3139 12484 3195 12486
rect 2899 11450 2955 11452
rect 2979 11450 3035 11452
rect 3059 11450 3115 11452
rect 3139 11450 3195 11452
rect 2899 11398 2945 11450
rect 2945 11398 2955 11450
rect 2979 11398 3009 11450
rect 3009 11398 3021 11450
rect 3021 11398 3035 11450
rect 3059 11398 3073 11450
rect 3073 11398 3085 11450
rect 3085 11398 3115 11450
rect 3139 11398 3149 11450
rect 3149 11398 3195 11450
rect 2899 11396 2955 11398
rect 2979 11396 3035 11398
rect 3059 11396 3115 11398
rect 3139 11396 3195 11398
rect 2899 10362 2955 10364
rect 2979 10362 3035 10364
rect 3059 10362 3115 10364
rect 3139 10362 3195 10364
rect 2899 10310 2945 10362
rect 2945 10310 2955 10362
rect 2979 10310 3009 10362
rect 3009 10310 3021 10362
rect 3021 10310 3035 10362
rect 3059 10310 3073 10362
rect 3073 10310 3085 10362
rect 3085 10310 3115 10362
rect 3139 10310 3149 10362
rect 3149 10310 3195 10362
rect 2899 10308 2955 10310
rect 2979 10308 3035 10310
rect 3059 10308 3115 10310
rect 3139 10308 3195 10310
rect 2899 9274 2955 9276
rect 2979 9274 3035 9276
rect 3059 9274 3115 9276
rect 3139 9274 3195 9276
rect 2899 9222 2945 9274
rect 2945 9222 2955 9274
rect 2979 9222 3009 9274
rect 3009 9222 3021 9274
rect 3021 9222 3035 9274
rect 3059 9222 3073 9274
rect 3073 9222 3085 9274
rect 3085 9222 3115 9274
rect 3139 9222 3149 9274
rect 3149 9222 3195 9274
rect 2899 9220 2955 9222
rect 2979 9220 3035 9222
rect 3059 9220 3115 9222
rect 3139 9220 3195 9222
rect 1398 8200 1454 8256
rect 2899 8186 2955 8188
rect 2979 8186 3035 8188
rect 3059 8186 3115 8188
rect 3139 8186 3195 8188
rect 2899 8134 2945 8186
rect 2945 8134 2955 8186
rect 2979 8134 3009 8186
rect 3009 8134 3021 8186
rect 3021 8134 3035 8186
rect 3059 8134 3073 8186
rect 3073 8134 3085 8186
rect 3085 8134 3115 8186
rect 3139 8134 3149 8186
rect 3149 8134 3195 8186
rect 2899 8132 2955 8134
rect 2979 8132 3035 8134
rect 3059 8132 3115 8134
rect 3139 8132 3195 8134
rect 4842 15258 4898 15260
rect 4922 15258 4978 15260
rect 5002 15258 5058 15260
rect 5082 15258 5138 15260
rect 4842 15206 4888 15258
rect 4888 15206 4898 15258
rect 4922 15206 4952 15258
rect 4952 15206 4964 15258
rect 4964 15206 4978 15258
rect 5002 15206 5016 15258
rect 5016 15206 5028 15258
rect 5028 15206 5058 15258
rect 5082 15206 5092 15258
rect 5092 15206 5138 15258
rect 4842 15204 4898 15206
rect 4922 15204 4978 15206
rect 5002 15204 5058 15206
rect 5082 15204 5138 15206
rect 4842 14170 4898 14172
rect 4922 14170 4978 14172
rect 5002 14170 5058 14172
rect 5082 14170 5138 14172
rect 4842 14118 4888 14170
rect 4888 14118 4898 14170
rect 4922 14118 4952 14170
rect 4952 14118 4964 14170
rect 4964 14118 4978 14170
rect 5002 14118 5016 14170
rect 5016 14118 5028 14170
rect 5028 14118 5058 14170
rect 5082 14118 5092 14170
rect 5092 14118 5138 14170
rect 4842 14116 4898 14118
rect 4922 14116 4978 14118
rect 5002 14116 5058 14118
rect 5082 14116 5138 14118
rect 2899 7098 2955 7100
rect 2979 7098 3035 7100
rect 3059 7098 3115 7100
rect 3139 7098 3195 7100
rect 2899 7046 2945 7098
rect 2945 7046 2955 7098
rect 2979 7046 3009 7098
rect 3009 7046 3021 7098
rect 3021 7046 3035 7098
rect 3059 7046 3073 7098
rect 3073 7046 3085 7098
rect 3085 7046 3115 7098
rect 3139 7046 3149 7098
rect 3149 7046 3195 7098
rect 2899 7044 2955 7046
rect 2979 7044 3035 7046
rect 3059 7044 3115 7046
rect 3139 7044 3195 7046
rect 2899 6010 2955 6012
rect 2979 6010 3035 6012
rect 3059 6010 3115 6012
rect 3139 6010 3195 6012
rect 2899 5958 2945 6010
rect 2945 5958 2955 6010
rect 2979 5958 3009 6010
rect 3009 5958 3021 6010
rect 3021 5958 3035 6010
rect 3059 5958 3073 6010
rect 3073 5958 3085 6010
rect 3085 5958 3115 6010
rect 3139 5958 3149 6010
rect 3149 5958 3195 6010
rect 2899 5956 2955 5958
rect 2979 5956 3035 5958
rect 3059 5956 3115 5958
rect 3139 5956 3195 5958
rect 4842 13082 4898 13084
rect 4922 13082 4978 13084
rect 5002 13082 5058 13084
rect 5082 13082 5138 13084
rect 4842 13030 4888 13082
rect 4888 13030 4898 13082
rect 4922 13030 4952 13082
rect 4952 13030 4964 13082
rect 4964 13030 4978 13082
rect 5002 13030 5016 13082
rect 5016 13030 5028 13082
rect 5028 13030 5058 13082
rect 5082 13030 5092 13082
rect 5092 13030 5138 13082
rect 4842 13028 4898 13030
rect 4922 13028 4978 13030
rect 5002 13028 5058 13030
rect 5082 13028 5138 13030
rect 5446 12688 5502 12744
rect 4842 11994 4898 11996
rect 4922 11994 4978 11996
rect 5002 11994 5058 11996
rect 5082 11994 5138 11996
rect 4842 11942 4888 11994
rect 4888 11942 4898 11994
rect 4922 11942 4952 11994
rect 4952 11942 4964 11994
rect 4964 11942 4978 11994
rect 5002 11942 5016 11994
rect 5016 11942 5028 11994
rect 5028 11942 5058 11994
rect 5082 11942 5092 11994
rect 5092 11942 5138 11994
rect 4842 11940 4898 11942
rect 4922 11940 4978 11942
rect 5002 11940 5058 11942
rect 5082 11940 5138 11942
rect 4842 10906 4898 10908
rect 4922 10906 4978 10908
rect 5002 10906 5058 10908
rect 5082 10906 5138 10908
rect 4842 10854 4888 10906
rect 4888 10854 4898 10906
rect 4922 10854 4952 10906
rect 4952 10854 4964 10906
rect 4964 10854 4978 10906
rect 5002 10854 5016 10906
rect 5016 10854 5028 10906
rect 5028 10854 5058 10906
rect 5082 10854 5092 10906
rect 5092 10854 5138 10906
rect 4842 10852 4898 10854
rect 4922 10852 4978 10854
rect 5002 10852 5058 10854
rect 5082 10852 5138 10854
rect 4842 9818 4898 9820
rect 4922 9818 4978 9820
rect 5002 9818 5058 9820
rect 5082 9818 5138 9820
rect 4842 9766 4888 9818
rect 4888 9766 4898 9818
rect 4922 9766 4952 9818
rect 4952 9766 4964 9818
rect 4964 9766 4978 9818
rect 5002 9766 5016 9818
rect 5016 9766 5028 9818
rect 5028 9766 5058 9818
rect 5082 9766 5092 9818
rect 5092 9766 5138 9818
rect 4842 9764 4898 9766
rect 4922 9764 4978 9766
rect 5002 9764 5058 9766
rect 5082 9764 5138 9766
rect 6786 15802 6842 15804
rect 6866 15802 6922 15804
rect 6946 15802 7002 15804
rect 7026 15802 7082 15804
rect 6786 15750 6832 15802
rect 6832 15750 6842 15802
rect 6866 15750 6896 15802
rect 6896 15750 6908 15802
rect 6908 15750 6922 15802
rect 6946 15750 6960 15802
rect 6960 15750 6972 15802
rect 6972 15750 7002 15802
rect 7026 15750 7036 15802
rect 7036 15750 7082 15802
rect 6786 15748 6842 15750
rect 6866 15748 6922 15750
rect 6946 15748 7002 15750
rect 7026 15748 7082 15750
rect 6786 14714 6842 14716
rect 6866 14714 6922 14716
rect 6946 14714 7002 14716
rect 7026 14714 7082 14716
rect 6786 14662 6832 14714
rect 6832 14662 6842 14714
rect 6866 14662 6896 14714
rect 6896 14662 6908 14714
rect 6908 14662 6922 14714
rect 6946 14662 6960 14714
rect 6960 14662 6972 14714
rect 6972 14662 7002 14714
rect 7026 14662 7036 14714
rect 7036 14662 7082 14714
rect 6786 14660 6842 14662
rect 6866 14660 6922 14662
rect 6946 14660 7002 14662
rect 7026 14660 7082 14662
rect 8729 16346 8785 16348
rect 8809 16346 8865 16348
rect 8889 16346 8945 16348
rect 8969 16346 9025 16348
rect 8729 16294 8775 16346
rect 8775 16294 8785 16346
rect 8809 16294 8839 16346
rect 8839 16294 8851 16346
rect 8851 16294 8865 16346
rect 8889 16294 8903 16346
rect 8903 16294 8915 16346
rect 8915 16294 8945 16346
rect 8969 16294 8979 16346
rect 8979 16294 9025 16346
rect 8729 16292 8785 16294
rect 8809 16292 8865 16294
rect 8889 16292 8945 16294
rect 8969 16292 9025 16294
rect 6786 13626 6842 13628
rect 6866 13626 6922 13628
rect 6946 13626 7002 13628
rect 7026 13626 7082 13628
rect 6786 13574 6832 13626
rect 6832 13574 6842 13626
rect 6866 13574 6896 13626
rect 6896 13574 6908 13626
rect 6908 13574 6922 13626
rect 6946 13574 6960 13626
rect 6960 13574 6972 13626
rect 6972 13574 7002 13626
rect 7026 13574 7036 13626
rect 7036 13574 7082 13626
rect 6786 13572 6842 13574
rect 6866 13572 6922 13574
rect 6946 13572 7002 13574
rect 7026 13572 7082 13574
rect 6786 12538 6842 12540
rect 6866 12538 6922 12540
rect 6946 12538 7002 12540
rect 7026 12538 7082 12540
rect 6786 12486 6832 12538
rect 6832 12486 6842 12538
rect 6866 12486 6896 12538
rect 6896 12486 6908 12538
rect 6908 12486 6922 12538
rect 6946 12486 6960 12538
rect 6960 12486 6972 12538
rect 6972 12486 7002 12538
rect 7026 12486 7036 12538
rect 7036 12486 7082 12538
rect 6786 12484 6842 12486
rect 6866 12484 6922 12486
rect 6946 12484 7002 12486
rect 7026 12484 7082 12486
rect 8729 15258 8785 15260
rect 8809 15258 8865 15260
rect 8889 15258 8945 15260
rect 8969 15258 9025 15260
rect 8729 15206 8775 15258
rect 8775 15206 8785 15258
rect 8809 15206 8839 15258
rect 8839 15206 8851 15258
rect 8851 15206 8865 15258
rect 8889 15206 8903 15258
rect 8903 15206 8915 15258
rect 8915 15206 8945 15258
rect 8969 15206 8979 15258
rect 8979 15206 9025 15258
rect 8729 15204 8785 15206
rect 8809 15204 8865 15206
rect 8889 15204 8945 15206
rect 8969 15204 9025 15206
rect 8729 14170 8785 14172
rect 8809 14170 8865 14172
rect 8889 14170 8945 14172
rect 8969 14170 9025 14172
rect 8729 14118 8775 14170
rect 8775 14118 8785 14170
rect 8809 14118 8839 14170
rect 8839 14118 8851 14170
rect 8851 14118 8865 14170
rect 8889 14118 8903 14170
rect 8903 14118 8915 14170
rect 8915 14118 8945 14170
rect 8969 14118 8979 14170
rect 8979 14118 9025 14170
rect 8729 14116 8785 14118
rect 8809 14116 8865 14118
rect 8889 14116 8945 14118
rect 8969 14116 9025 14118
rect 8729 13082 8785 13084
rect 8809 13082 8865 13084
rect 8889 13082 8945 13084
rect 8969 13082 9025 13084
rect 8729 13030 8775 13082
rect 8775 13030 8785 13082
rect 8809 13030 8839 13082
rect 8839 13030 8851 13082
rect 8851 13030 8865 13082
rect 8889 13030 8903 13082
rect 8903 13030 8915 13082
rect 8915 13030 8945 13082
rect 8969 13030 8979 13082
rect 8979 13030 9025 13082
rect 8729 13028 8785 13030
rect 8809 13028 8865 13030
rect 8889 13028 8945 13030
rect 8969 13028 9025 13030
rect 6786 11450 6842 11452
rect 6866 11450 6922 11452
rect 6946 11450 7002 11452
rect 7026 11450 7082 11452
rect 6786 11398 6832 11450
rect 6832 11398 6842 11450
rect 6866 11398 6896 11450
rect 6896 11398 6908 11450
rect 6908 11398 6922 11450
rect 6946 11398 6960 11450
rect 6960 11398 6972 11450
rect 6972 11398 7002 11450
rect 7026 11398 7036 11450
rect 7036 11398 7082 11450
rect 6786 11396 6842 11398
rect 6866 11396 6922 11398
rect 6946 11396 7002 11398
rect 7026 11396 7082 11398
rect 6786 10362 6842 10364
rect 6866 10362 6922 10364
rect 6946 10362 7002 10364
rect 7026 10362 7082 10364
rect 6786 10310 6832 10362
rect 6832 10310 6842 10362
rect 6866 10310 6896 10362
rect 6896 10310 6908 10362
rect 6908 10310 6922 10362
rect 6946 10310 6960 10362
rect 6960 10310 6972 10362
rect 6972 10310 7002 10362
rect 7026 10310 7036 10362
rect 7036 10310 7082 10362
rect 6786 10308 6842 10310
rect 6866 10308 6922 10310
rect 6946 10308 7002 10310
rect 7026 10308 7082 10310
rect 4842 8730 4898 8732
rect 4922 8730 4978 8732
rect 5002 8730 5058 8732
rect 5082 8730 5138 8732
rect 4842 8678 4888 8730
rect 4888 8678 4898 8730
rect 4922 8678 4952 8730
rect 4952 8678 4964 8730
rect 4964 8678 4978 8730
rect 5002 8678 5016 8730
rect 5016 8678 5028 8730
rect 5028 8678 5058 8730
rect 5082 8678 5092 8730
rect 5092 8678 5138 8730
rect 4842 8676 4898 8678
rect 4922 8676 4978 8678
rect 5002 8676 5058 8678
rect 5082 8676 5138 8678
rect 938 4156 940 4176
rect 940 4156 992 4176
rect 992 4156 994 4176
rect 938 4120 994 4156
rect 2899 4922 2955 4924
rect 2979 4922 3035 4924
rect 3059 4922 3115 4924
rect 3139 4922 3195 4924
rect 2899 4870 2945 4922
rect 2945 4870 2955 4922
rect 2979 4870 3009 4922
rect 3009 4870 3021 4922
rect 3021 4870 3035 4922
rect 3059 4870 3073 4922
rect 3073 4870 3085 4922
rect 3085 4870 3115 4922
rect 3139 4870 3149 4922
rect 3149 4870 3195 4922
rect 2899 4868 2955 4870
rect 2979 4868 3035 4870
rect 3059 4868 3115 4870
rect 3139 4868 3195 4870
rect 2899 3834 2955 3836
rect 2979 3834 3035 3836
rect 3059 3834 3115 3836
rect 3139 3834 3195 3836
rect 2899 3782 2945 3834
rect 2945 3782 2955 3834
rect 2979 3782 3009 3834
rect 3009 3782 3021 3834
rect 3021 3782 3035 3834
rect 3059 3782 3073 3834
rect 3073 3782 3085 3834
rect 3085 3782 3115 3834
rect 3139 3782 3149 3834
rect 3149 3782 3195 3834
rect 2899 3780 2955 3782
rect 2979 3780 3035 3782
rect 3059 3780 3115 3782
rect 3139 3780 3195 3782
rect 2899 2746 2955 2748
rect 2979 2746 3035 2748
rect 3059 2746 3115 2748
rect 3139 2746 3195 2748
rect 2899 2694 2945 2746
rect 2945 2694 2955 2746
rect 2979 2694 3009 2746
rect 3009 2694 3021 2746
rect 3021 2694 3035 2746
rect 3059 2694 3073 2746
rect 3073 2694 3085 2746
rect 3085 2694 3115 2746
rect 3139 2694 3149 2746
rect 3149 2694 3195 2746
rect 2899 2692 2955 2694
rect 2979 2692 3035 2694
rect 3059 2692 3115 2694
rect 3139 2692 3195 2694
rect 4842 7642 4898 7644
rect 4922 7642 4978 7644
rect 5002 7642 5058 7644
rect 5082 7642 5138 7644
rect 4842 7590 4888 7642
rect 4888 7590 4898 7642
rect 4922 7590 4952 7642
rect 4952 7590 4964 7642
rect 4964 7590 4978 7642
rect 5002 7590 5016 7642
rect 5016 7590 5028 7642
rect 5028 7590 5058 7642
rect 5082 7590 5092 7642
rect 5092 7590 5138 7642
rect 4842 7588 4898 7590
rect 4922 7588 4978 7590
rect 5002 7588 5058 7590
rect 5082 7588 5138 7590
rect 4842 6554 4898 6556
rect 4922 6554 4978 6556
rect 5002 6554 5058 6556
rect 5082 6554 5138 6556
rect 4842 6502 4888 6554
rect 4888 6502 4898 6554
rect 4922 6502 4952 6554
rect 4952 6502 4964 6554
rect 4964 6502 4978 6554
rect 5002 6502 5016 6554
rect 5016 6502 5028 6554
rect 5028 6502 5058 6554
rect 5082 6502 5092 6554
rect 5092 6502 5138 6554
rect 4842 6500 4898 6502
rect 4922 6500 4978 6502
rect 5002 6500 5058 6502
rect 5082 6500 5138 6502
rect 4842 5466 4898 5468
rect 4922 5466 4978 5468
rect 5002 5466 5058 5468
rect 5082 5466 5138 5468
rect 4842 5414 4888 5466
rect 4888 5414 4898 5466
rect 4922 5414 4952 5466
rect 4952 5414 4964 5466
rect 4964 5414 4978 5466
rect 5002 5414 5016 5466
rect 5016 5414 5028 5466
rect 5028 5414 5058 5466
rect 5082 5414 5092 5466
rect 5092 5414 5138 5466
rect 4842 5412 4898 5414
rect 4922 5412 4978 5414
rect 5002 5412 5058 5414
rect 5082 5412 5138 5414
rect 6786 9274 6842 9276
rect 6866 9274 6922 9276
rect 6946 9274 7002 9276
rect 7026 9274 7082 9276
rect 6786 9222 6832 9274
rect 6832 9222 6842 9274
rect 6866 9222 6896 9274
rect 6896 9222 6908 9274
rect 6908 9222 6922 9274
rect 6946 9222 6960 9274
rect 6960 9222 6972 9274
rect 6972 9222 7002 9274
rect 7026 9222 7036 9274
rect 7036 9222 7082 9274
rect 6786 9220 6842 9222
rect 6866 9220 6922 9222
rect 6946 9220 7002 9222
rect 7026 9220 7082 9222
rect 8729 11994 8785 11996
rect 8809 11994 8865 11996
rect 8889 11994 8945 11996
rect 8969 11994 9025 11996
rect 8729 11942 8775 11994
rect 8775 11942 8785 11994
rect 8809 11942 8839 11994
rect 8839 11942 8851 11994
rect 8851 11942 8865 11994
rect 8889 11942 8903 11994
rect 8903 11942 8915 11994
rect 8915 11942 8945 11994
rect 8969 11942 8979 11994
rect 8979 11942 9025 11994
rect 8729 11940 8785 11942
rect 8809 11940 8865 11942
rect 8889 11940 8945 11942
rect 8969 11940 9025 11942
rect 8729 10906 8785 10908
rect 8809 10906 8865 10908
rect 8889 10906 8945 10908
rect 8969 10906 9025 10908
rect 8729 10854 8775 10906
rect 8775 10854 8785 10906
rect 8809 10854 8839 10906
rect 8839 10854 8851 10906
rect 8851 10854 8865 10906
rect 8889 10854 8903 10906
rect 8903 10854 8915 10906
rect 8915 10854 8945 10906
rect 8969 10854 8979 10906
rect 8979 10854 9025 10906
rect 8729 10852 8785 10854
rect 8809 10852 8865 10854
rect 8889 10852 8945 10854
rect 8969 10852 9025 10854
rect 6786 8186 6842 8188
rect 6866 8186 6922 8188
rect 6946 8186 7002 8188
rect 7026 8186 7082 8188
rect 6786 8134 6832 8186
rect 6832 8134 6842 8186
rect 6866 8134 6896 8186
rect 6896 8134 6908 8186
rect 6908 8134 6922 8186
rect 6946 8134 6960 8186
rect 6960 8134 6972 8186
rect 6972 8134 7002 8186
rect 7026 8134 7036 8186
rect 7036 8134 7082 8186
rect 6786 8132 6842 8134
rect 6866 8132 6922 8134
rect 6946 8132 7002 8134
rect 7026 8132 7082 8134
rect 6786 7098 6842 7100
rect 6866 7098 6922 7100
rect 6946 7098 7002 7100
rect 7026 7098 7082 7100
rect 6786 7046 6832 7098
rect 6832 7046 6842 7098
rect 6866 7046 6896 7098
rect 6896 7046 6908 7098
rect 6908 7046 6922 7098
rect 6946 7046 6960 7098
rect 6960 7046 6972 7098
rect 6972 7046 7002 7098
rect 7026 7046 7036 7098
rect 7036 7046 7082 7098
rect 6786 7044 6842 7046
rect 6866 7044 6922 7046
rect 6946 7044 7002 7046
rect 7026 7044 7082 7046
rect 4842 4378 4898 4380
rect 4922 4378 4978 4380
rect 5002 4378 5058 4380
rect 5082 4378 5138 4380
rect 4842 4326 4888 4378
rect 4888 4326 4898 4378
rect 4922 4326 4952 4378
rect 4952 4326 4964 4378
rect 4964 4326 4978 4378
rect 5002 4326 5016 4378
rect 5016 4326 5028 4378
rect 5028 4326 5058 4378
rect 5082 4326 5092 4378
rect 5092 4326 5138 4378
rect 4842 4324 4898 4326
rect 4922 4324 4978 4326
rect 5002 4324 5058 4326
rect 5082 4324 5138 4326
rect 4842 3290 4898 3292
rect 4922 3290 4978 3292
rect 5002 3290 5058 3292
rect 5082 3290 5138 3292
rect 4842 3238 4888 3290
rect 4888 3238 4898 3290
rect 4922 3238 4952 3290
rect 4952 3238 4964 3290
rect 4964 3238 4978 3290
rect 5002 3238 5016 3290
rect 5016 3238 5028 3290
rect 5028 3238 5058 3290
rect 5082 3238 5092 3290
rect 5092 3238 5138 3290
rect 4842 3236 4898 3238
rect 4922 3236 4978 3238
rect 5002 3236 5058 3238
rect 5082 3236 5138 3238
rect 6786 6010 6842 6012
rect 6866 6010 6922 6012
rect 6946 6010 7002 6012
rect 7026 6010 7082 6012
rect 6786 5958 6832 6010
rect 6832 5958 6842 6010
rect 6866 5958 6896 6010
rect 6896 5958 6908 6010
rect 6908 5958 6922 6010
rect 6946 5958 6960 6010
rect 6960 5958 6972 6010
rect 6972 5958 7002 6010
rect 7026 5958 7036 6010
rect 7036 5958 7082 6010
rect 6786 5956 6842 5958
rect 6866 5956 6922 5958
rect 6946 5956 7002 5958
rect 7026 5956 7082 5958
rect 6786 4922 6842 4924
rect 6866 4922 6922 4924
rect 6946 4922 7002 4924
rect 7026 4922 7082 4924
rect 6786 4870 6832 4922
rect 6832 4870 6842 4922
rect 6866 4870 6896 4922
rect 6896 4870 6908 4922
rect 6908 4870 6922 4922
rect 6946 4870 6960 4922
rect 6960 4870 6972 4922
rect 6972 4870 7002 4922
rect 7026 4870 7036 4922
rect 7036 4870 7082 4922
rect 6786 4868 6842 4870
rect 6866 4868 6922 4870
rect 6946 4868 7002 4870
rect 7026 4868 7082 4870
rect 6786 3834 6842 3836
rect 6866 3834 6922 3836
rect 6946 3834 7002 3836
rect 7026 3834 7082 3836
rect 6786 3782 6832 3834
rect 6832 3782 6842 3834
rect 6866 3782 6896 3834
rect 6896 3782 6908 3834
rect 6908 3782 6922 3834
rect 6946 3782 6960 3834
rect 6960 3782 6972 3834
rect 6972 3782 7002 3834
rect 7026 3782 7036 3834
rect 7036 3782 7082 3834
rect 6786 3780 6842 3782
rect 6866 3780 6922 3782
rect 6946 3780 7002 3782
rect 7026 3780 7082 3782
rect 6786 2746 6842 2748
rect 6866 2746 6922 2748
rect 6946 2746 7002 2748
rect 7026 2746 7082 2748
rect 6786 2694 6832 2746
rect 6832 2694 6842 2746
rect 6866 2694 6896 2746
rect 6896 2694 6908 2746
rect 6908 2694 6922 2746
rect 6946 2694 6960 2746
rect 6960 2694 6972 2746
rect 6972 2694 7002 2746
rect 7026 2694 7036 2746
rect 7036 2694 7082 2746
rect 6786 2692 6842 2694
rect 6866 2692 6922 2694
rect 6946 2692 7002 2694
rect 7026 2692 7082 2694
rect 8729 9818 8785 9820
rect 8809 9818 8865 9820
rect 8889 9818 8945 9820
rect 8969 9818 9025 9820
rect 8729 9766 8775 9818
rect 8775 9766 8785 9818
rect 8809 9766 8839 9818
rect 8839 9766 8851 9818
rect 8851 9766 8865 9818
rect 8889 9766 8903 9818
rect 8903 9766 8915 9818
rect 8915 9766 8945 9818
rect 8969 9766 8979 9818
rect 8979 9766 9025 9818
rect 8729 9764 8785 9766
rect 8809 9764 8865 9766
rect 8889 9764 8945 9766
rect 8969 9764 9025 9766
rect 8729 8730 8785 8732
rect 8809 8730 8865 8732
rect 8889 8730 8945 8732
rect 8969 8730 9025 8732
rect 8729 8678 8775 8730
rect 8775 8678 8785 8730
rect 8809 8678 8839 8730
rect 8839 8678 8851 8730
rect 8851 8678 8865 8730
rect 8889 8678 8903 8730
rect 8903 8678 8915 8730
rect 8915 8678 8945 8730
rect 8969 8678 8979 8730
rect 8979 8678 9025 8730
rect 8729 8676 8785 8678
rect 8809 8676 8865 8678
rect 8889 8676 8945 8678
rect 8969 8676 9025 8678
rect 9862 12688 9918 12744
rect 8729 7642 8785 7644
rect 8809 7642 8865 7644
rect 8889 7642 8945 7644
rect 8969 7642 9025 7644
rect 8729 7590 8775 7642
rect 8775 7590 8785 7642
rect 8809 7590 8839 7642
rect 8839 7590 8851 7642
rect 8851 7590 8865 7642
rect 8889 7590 8903 7642
rect 8903 7590 8915 7642
rect 8915 7590 8945 7642
rect 8969 7590 8979 7642
rect 8979 7590 9025 7642
rect 8729 7588 8785 7590
rect 8809 7588 8865 7590
rect 8889 7588 8945 7590
rect 8969 7588 9025 7590
rect 8729 6554 8785 6556
rect 8809 6554 8865 6556
rect 8889 6554 8945 6556
rect 8969 6554 9025 6556
rect 8729 6502 8775 6554
rect 8775 6502 8785 6554
rect 8809 6502 8839 6554
rect 8839 6502 8851 6554
rect 8851 6502 8865 6554
rect 8889 6502 8903 6554
rect 8903 6502 8915 6554
rect 8915 6502 8945 6554
rect 8969 6502 8979 6554
rect 8979 6502 9025 6554
rect 8729 6500 8785 6502
rect 8809 6500 8865 6502
rect 8889 6500 8945 6502
rect 8969 6500 9025 6502
rect 8729 5466 8785 5468
rect 8809 5466 8865 5468
rect 8889 5466 8945 5468
rect 8969 5466 9025 5468
rect 8729 5414 8775 5466
rect 8775 5414 8785 5466
rect 8809 5414 8839 5466
rect 8839 5414 8851 5466
rect 8851 5414 8865 5466
rect 8889 5414 8903 5466
rect 8903 5414 8915 5466
rect 8915 5414 8945 5466
rect 8969 5414 8979 5466
rect 8979 5414 9025 5466
rect 8729 5412 8785 5414
rect 8809 5412 8865 5414
rect 8889 5412 8945 5414
rect 8969 5412 9025 5414
rect 8729 4378 8785 4380
rect 8809 4378 8865 4380
rect 8889 4378 8945 4380
rect 8969 4378 9025 4380
rect 8729 4326 8775 4378
rect 8775 4326 8785 4378
rect 8809 4326 8839 4378
rect 8839 4326 8851 4378
rect 8851 4326 8865 4378
rect 8889 4326 8903 4378
rect 8903 4326 8915 4378
rect 8915 4326 8945 4378
rect 8969 4326 8979 4378
rect 8979 4326 9025 4378
rect 8729 4324 8785 4326
rect 8809 4324 8865 4326
rect 8889 4324 8945 4326
rect 8969 4324 9025 4326
rect 8729 3290 8785 3292
rect 8809 3290 8865 3292
rect 8889 3290 8945 3292
rect 8969 3290 9025 3292
rect 8729 3238 8775 3290
rect 8775 3238 8785 3290
rect 8809 3238 8839 3290
rect 8839 3238 8851 3290
rect 8851 3238 8865 3290
rect 8889 3238 8903 3290
rect 8903 3238 8915 3290
rect 8915 3238 8945 3290
rect 8969 3238 8979 3290
rect 8979 3238 9025 3290
rect 8729 3236 8785 3238
rect 8809 3236 8865 3238
rect 8889 3236 8945 3238
rect 8969 3236 9025 3238
rect 10673 16890 10729 16892
rect 10753 16890 10809 16892
rect 10833 16890 10889 16892
rect 10913 16890 10969 16892
rect 10673 16838 10719 16890
rect 10719 16838 10729 16890
rect 10753 16838 10783 16890
rect 10783 16838 10795 16890
rect 10795 16838 10809 16890
rect 10833 16838 10847 16890
rect 10847 16838 10859 16890
rect 10859 16838 10889 16890
rect 10913 16838 10923 16890
rect 10923 16838 10969 16890
rect 10673 16836 10729 16838
rect 10753 16836 10809 16838
rect 10833 16836 10889 16838
rect 10913 16836 10969 16838
rect 10673 15802 10729 15804
rect 10753 15802 10809 15804
rect 10833 15802 10889 15804
rect 10913 15802 10969 15804
rect 10673 15750 10719 15802
rect 10719 15750 10729 15802
rect 10753 15750 10783 15802
rect 10783 15750 10795 15802
rect 10795 15750 10809 15802
rect 10833 15750 10847 15802
rect 10847 15750 10859 15802
rect 10859 15750 10889 15802
rect 10913 15750 10923 15802
rect 10923 15750 10969 15802
rect 10673 15748 10729 15750
rect 10753 15748 10809 15750
rect 10833 15748 10889 15750
rect 10913 15748 10969 15750
rect 10673 14714 10729 14716
rect 10753 14714 10809 14716
rect 10833 14714 10889 14716
rect 10913 14714 10969 14716
rect 10673 14662 10719 14714
rect 10719 14662 10729 14714
rect 10753 14662 10783 14714
rect 10783 14662 10795 14714
rect 10795 14662 10809 14714
rect 10833 14662 10847 14714
rect 10847 14662 10859 14714
rect 10859 14662 10889 14714
rect 10913 14662 10923 14714
rect 10923 14662 10969 14714
rect 10673 14660 10729 14662
rect 10753 14660 10809 14662
rect 10833 14660 10889 14662
rect 10913 14660 10969 14662
rect 14560 16890 14616 16892
rect 14640 16890 14696 16892
rect 14720 16890 14776 16892
rect 14800 16890 14856 16892
rect 14560 16838 14606 16890
rect 14606 16838 14616 16890
rect 14640 16838 14670 16890
rect 14670 16838 14682 16890
rect 14682 16838 14696 16890
rect 14720 16838 14734 16890
rect 14734 16838 14746 16890
rect 14746 16838 14776 16890
rect 14800 16838 14810 16890
rect 14810 16838 14856 16890
rect 14560 16836 14616 16838
rect 14640 16836 14696 16838
rect 14720 16836 14776 16838
rect 14800 16836 14856 16838
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 10673 13626 10729 13628
rect 10753 13626 10809 13628
rect 10833 13626 10889 13628
rect 10913 13626 10969 13628
rect 10673 13574 10719 13626
rect 10719 13574 10729 13626
rect 10753 13574 10783 13626
rect 10783 13574 10795 13626
rect 10795 13574 10809 13626
rect 10833 13574 10847 13626
rect 10847 13574 10859 13626
rect 10859 13574 10889 13626
rect 10913 13574 10923 13626
rect 10923 13574 10969 13626
rect 10673 13572 10729 13574
rect 10753 13572 10809 13574
rect 10833 13572 10889 13574
rect 10913 13572 10969 13574
rect 10673 12538 10729 12540
rect 10753 12538 10809 12540
rect 10833 12538 10889 12540
rect 10913 12538 10969 12540
rect 10673 12486 10719 12538
rect 10719 12486 10729 12538
rect 10753 12486 10783 12538
rect 10783 12486 10795 12538
rect 10795 12486 10809 12538
rect 10833 12486 10847 12538
rect 10847 12486 10859 12538
rect 10859 12486 10889 12538
rect 10913 12486 10923 12538
rect 10923 12486 10969 12538
rect 10673 12484 10729 12486
rect 10753 12484 10809 12486
rect 10833 12484 10889 12486
rect 10913 12484 10969 12486
rect 10673 11450 10729 11452
rect 10753 11450 10809 11452
rect 10833 11450 10889 11452
rect 10913 11450 10969 11452
rect 10673 11398 10719 11450
rect 10719 11398 10729 11450
rect 10753 11398 10783 11450
rect 10783 11398 10795 11450
rect 10795 11398 10809 11450
rect 10833 11398 10847 11450
rect 10847 11398 10859 11450
rect 10859 11398 10889 11450
rect 10913 11398 10923 11450
rect 10923 11398 10969 11450
rect 10673 11396 10729 11398
rect 10753 11396 10809 11398
rect 10833 11396 10889 11398
rect 10913 11396 10969 11398
rect 10673 10362 10729 10364
rect 10753 10362 10809 10364
rect 10833 10362 10889 10364
rect 10913 10362 10969 10364
rect 10673 10310 10719 10362
rect 10719 10310 10729 10362
rect 10753 10310 10783 10362
rect 10783 10310 10795 10362
rect 10795 10310 10809 10362
rect 10833 10310 10847 10362
rect 10847 10310 10859 10362
rect 10859 10310 10889 10362
rect 10913 10310 10923 10362
rect 10923 10310 10969 10362
rect 10673 10308 10729 10310
rect 10753 10308 10809 10310
rect 10833 10308 10889 10310
rect 10913 10308 10969 10310
rect 10673 9274 10729 9276
rect 10753 9274 10809 9276
rect 10833 9274 10889 9276
rect 10913 9274 10969 9276
rect 10673 9222 10719 9274
rect 10719 9222 10729 9274
rect 10753 9222 10783 9274
rect 10783 9222 10795 9274
rect 10795 9222 10809 9274
rect 10833 9222 10847 9274
rect 10847 9222 10859 9274
rect 10859 9222 10889 9274
rect 10913 9222 10923 9274
rect 10923 9222 10969 9274
rect 10673 9220 10729 9222
rect 10753 9220 10809 9222
rect 10833 9220 10889 9222
rect 10913 9220 10969 9222
rect 10673 8186 10729 8188
rect 10753 8186 10809 8188
rect 10833 8186 10889 8188
rect 10913 8186 10969 8188
rect 10673 8134 10719 8186
rect 10719 8134 10729 8186
rect 10753 8134 10783 8186
rect 10783 8134 10795 8186
rect 10795 8134 10809 8186
rect 10833 8134 10847 8186
rect 10847 8134 10859 8186
rect 10859 8134 10889 8186
rect 10913 8134 10923 8186
rect 10923 8134 10969 8186
rect 10673 8132 10729 8134
rect 10753 8132 10809 8134
rect 10833 8132 10889 8134
rect 10913 8132 10969 8134
rect 10673 7098 10729 7100
rect 10753 7098 10809 7100
rect 10833 7098 10889 7100
rect 10913 7098 10969 7100
rect 10673 7046 10719 7098
rect 10719 7046 10729 7098
rect 10753 7046 10783 7098
rect 10783 7046 10795 7098
rect 10795 7046 10809 7098
rect 10833 7046 10847 7098
rect 10847 7046 10859 7098
rect 10859 7046 10889 7098
rect 10913 7046 10923 7098
rect 10923 7046 10969 7098
rect 10673 7044 10729 7046
rect 10753 7044 10809 7046
rect 10833 7044 10889 7046
rect 10913 7044 10969 7046
rect 10673 6010 10729 6012
rect 10753 6010 10809 6012
rect 10833 6010 10889 6012
rect 10913 6010 10969 6012
rect 10673 5958 10719 6010
rect 10719 5958 10729 6010
rect 10753 5958 10783 6010
rect 10783 5958 10795 6010
rect 10795 5958 10809 6010
rect 10833 5958 10847 6010
rect 10847 5958 10859 6010
rect 10859 5958 10889 6010
rect 10913 5958 10923 6010
rect 10923 5958 10969 6010
rect 10673 5956 10729 5958
rect 10753 5956 10809 5958
rect 10833 5956 10889 5958
rect 10913 5956 10969 5958
rect 14560 15802 14616 15804
rect 14640 15802 14696 15804
rect 14720 15802 14776 15804
rect 14800 15802 14856 15804
rect 14560 15750 14606 15802
rect 14606 15750 14616 15802
rect 14640 15750 14670 15802
rect 14670 15750 14682 15802
rect 14682 15750 14696 15802
rect 14720 15750 14734 15802
rect 14734 15750 14746 15802
rect 14746 15750 14776 15802
rect 14800 15750 14810 15802
rect 14810 15750 14856 15802
rect 14560 15748 14616 15750
rect 14640 15748 14696 15750
rect 14720 15748 14776 15750
rect 14800 15748 14856 15750
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 14560 14714 14616 14716
rect 14640 14714 14696 14716
rect 14720 14714 14776 14716
rect 14800 14714 14856 14716
rect 14560 14662 14606 14714
rect 14606 14662 14616 14714
rect 14640 14662 14670 14714
rect 14670 14662 14682 14714
rect 14682 14662 14696 14714
rect 14720 14662 14734 14714
rect 14734 14662 14746 14714
rect 14746 14662 14776 14714
rect 14800 14662 14810 14714
rect 14810 14662 14856 14714
rect 14560 14660 14616 14662
rect 14640 14660 14696 14662
rect 14720 14660 14776 14662
rect 14800 14660 14856 14662
rect 14560 13626 14616 13628
rect 14640 13626 14696 13628
rect 14720 13626 14776 13628
rect 14800 13626 14856 13628
rect 14560 13574 14606 13626
rect 14606 13574 14616 13626
rect 14640 13574 14670 13626
rect 14670 13574 14682 13626
rect 14682 13574 14696 13626
rect 14720 13574 14734 13626
rect 14734 13574 14746 13626
rect 14746 13574 14776 13626
rect 14800 13574 14810 13626
rect 14810 13574 14856 13626
rect 14560 13572 14616 13574
rect 14640 13572 14696 13574
rect 14720 13572 14776 13574
rect 14800 13572 14856 13574
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 14560 12538 14616 12540
rect 14640 12538 14696 12540
rect 14720 12538 14776 12540
rect 14800 12538 14856 12540
rect 14560 12486 14606 12538
rect 14606 12486 14616 12538
rect 14640 12486 14670 12538
rect 14670 12486 14682 12538
rect 14682 12486 14696 12538
rect 14720 12486 14734 12538
rect 14734 12486 14746 12538
rect 14746 12486 14776 12538
rect 14800 12486 14810 12538
rect 14810 12486 14856 12538
rect 14560 12484 14616 12486
rect 14640 12484 14696 12486
rect 14720 12484 14776 12486
rect 14800 12484 14856 12486
rect 16503 16346 16559 16348
rect 16583 16346 16639 16348
rect 16663 16346 16719 16348
rect 16743 16346 16799 16348
rect 16503 16294 16549 16346
rect 16549 16294 16559 16346
rect 16583 16294 16613 16346
rect 16613 16294 16625 16346
rect 16625 16294 16639 16346
rect 16663 16294 16677 16346
rect 16677 16294 16689 16346
rect 16689 16294 16719 16346
rect 16743 16294 16753 16346
rect 16753 16294 16799 16346
rect 16503 16292 16559 16294
rect 16583 16292 16639 16294
rect 16663 16292 16719 16294
rect 16743 16292 16799 16294
rect 16503 15258 16559 15260
rect 16583 15258 16639 15260
rect 16663 15258 16719 15260
rect 16743 15258 16799 15260
rect 16503 15206 16549 15258
rect 16549 15206 16559 15258
rect 16583 15206 16613 15258
rect 16613 15206 16625 15258
rect 16625 15206 16639 15258
rect 16663 15206 16677 15258
rect 16677 15206 16689 15258
rect 16689 15206 16719 15258
rect 16743 15206 16753 15258
rect 16753 15206 16799 15258
rect 16503 15204 16559 15206
rect 16583 15204 16639 15206
rect 16663 15204 16719 15206
rect 16743 15204 16799 15206
rect 16503 14170 16559 14172
rect 16583 14170 16639 14172
rect 16663 14170 16719 14172
rect 16743 14170 16799 14172
rect 16503 14118 16549 14170
rect 16549 14118 16559 14170
rect 16583 14118 16613 14170
rect 16613 14118 16625 14170
rect 16625 14118 16639 14170
rect 16663 14118 16677 14170
rect 16677 14118 16689 14170
rect 16689 14118 16719 14170
rect 16743 14118 16753 14170
rect 16753 14118 16799 14170
rect 16503 14116 16559 14118
rect 16583 14116 16639 14118
rect 16663 14116 16719 14118
rect 16743 14116 16799 14118
rect 16578 13640 16634 13696
rect 16503 13082 16559 13084
rect 16583 13082 16639 13084
rect 16663 13082 16719 13084
rect 16743 13082 16799 13084
rect 16503 13030 16549 13082
rect 16549 13030 16559 13082
rect 16583 13030 16613 13082
rect 16613 13030 16625 13082
rect 16625 13030 16639 13082
rect 16663 13030 16677 13082
rect 16677 13030 16689 13082
rect 16689 13030 16719 13082
rect 16743 13030 16753 13082
rect 16753 13030 16799 13082
rect 16503 13028 16559 13030
rect 16583 13028 16639 13030
rect 16663 13028 16719 13030
rect 16743 13028 16799 13030
rect 14560 11450 14616 11452
rect 14640 11450 14696 11452
rect 14720 11450 14776 11452
rect 14800 11450 14856 11452
rect 14560 11398 14606 11450
rect 14606 11398 14616 11450
rect 14640 11398 14670 11450
rect 14670 11398 14682 11450
rect 14682 11398 14696 11450
rect 14720 11398 14734 11450
rect 14734 11398 14746 11450
rect 14746 11398 14776 11450
rect 14800 11398 14810 11450
rect 14810 11398 14856 11450
rect 14560 11396 14616 11398
rect 14640 11396 14696 11398
rect 14720 11396 14776 11398
rect 14800 11396 14856 11398
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 10673 4922 10729 4924
rect 10753 4922 10809 4924
rect 10833 4922 10889 4924
rect 10913 4922 10969 4924
rect 10673 4870 10719 4922
rect 10719 4870 10729 4922
rect 10753 4870 10783 4922
rect 10783 4870 10795 4922
rect 10795 4870 10809 4922
rect 10833 4870 10847 4922
rect 10847 4870 10859 4922
rect 10859 4870 10889 4922
rect 10913 4870 10923 4922
rect 10923 4870 10969 4922
rect 10673 4868 10729 4870
rect 10753 4868 10809 4870
rect 10833 4868 10889 4870
rect 10913 4868 10969 4870
rect 10673 3834 10729 3836
rect 10753 3834 10809 3836
rect 10833 3834 10889 3836
rect 10913 3834 10969 3836
rect 10673 3782 10719 3834
rect 10719 3782 10729 3834
rect 10753 3782 10783 3834
rect 10783 3782 10795 3834
rect 10795 3782 10809 3834
rect 10833 3782 10847 3834
rect 10847 3782 10859 3834
rect 10859 3782 10889 3834
rect 10913 3782 10923 3834
rect 10923 3782 10969 3834
rect 10673 3780 10729 3782
rect 10753 3780 10809 3782
rect 10833 3780 10889 3782
rect 10913 3780 10969 3782
rect 4842 2202 4898 2204
rect 4922 2202 4978 2204
rect 5002 2202 5058 2204
rect 5082 2202 5138 2204
rect 4842 2150 4888 2202
rect 4888 2150 4898 2202
rect 4922 2150 4952 2202
rect 4952 2150 4964 2202
rect 4964 2150 4978 2202
rect 5002 2150 5016 2202
rect 5016 2150 5028 2202
rect 5028 2150 5058 2202
rect 5082 2150 5092 2202
rect 5092 2150 5138 2202
rect 4842 2148 4898 2150
rect 4922 2148 4978 2150
rect 5002 2148 5058 2150
rect 5082 2148 5138 2150
rect 10673 2746 10729 2748
rect 10753 2746 10809 2748
rect 10833 2746 10889 2748
rect 10913 2746 10969 2748
rect 10673 2694 10719 2746
rect 10719 2694 10729 2746
rect 10753 2694 10783 2746
rect 10783 2694 10795 2746
rect 10795 2694 10809 2746
rect 10833 2694 10847 2746
rect 10847 2694 10859 2746
rect 10859 2694 10889 2746
rect 10913 2694 10923 2746
rect 10923 2694 10969 2746
rect 10673 2692 10729 2694
rect 10753 2692 10809 2694
rect 10833 2692 10889 2694
rect 10913 2692 10969 2694
rect 8729 2202 8785 2204
rect 8809 2202 8865 2204
rect 8889 2202 8945 2204
rect 8969 2202 9025 2204
rect 8729 2150 8775 2202
rect 8775 2150 8785 2202
rect 8809 2150 8839 2202
rect 8839 2150 8851 2202
rect 8851 2150 8865 2202
rect 8889 2150 8903 2202
rect 8903 2150 8915 2202
rect 8915 2150 8945 2202
rect 8969 2150 8979 2202
rect 8979 2150 9025 2202
rect 8729 2148 8785 2150
rect 8809 2148 8865 2150
rect 8889 2148 8945 2150
rect 8969 2148 9025 2150
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 14560 10362 14616 10364
rect 14640 10362 14696 10364
rect 14720 10362 14776 10364
rect 14800 10362 14856 10364
rect 14560 10310 14606 10362
rect 14606 10310 14616 10362
rect 14640 10310 14670 10362
rect 14670 10310 14682 10362
rect 14682 10310 14696 10362
rect 14720 10310 14734 10362
rect 14734 10310 14746 10362
rect 14746 10310 14776 10362
rect 14800 10310 14810 10362
rect 14810 10310 14856 10362
rect 14560 10308 14616 10310
rect 14640 10308 14696 10310
rect 14720 10308 14776 10310
rect 14800 10308 14856 10310
rect 16503 11994 16559 11996
rect 16583 11994 16639 11996
rect 16663 11994 16719 11996
rect 16743 11994 16799 11996
rect 16503 11942 16549 11994
rect 16549 11942 16559 11994
rect 16583 11942 16613 11994
rect 16613 11942 16625 11994
rect 16625 11942 16639 11994
rect 16663 11942 16677 11994
rect 16677 11942 16689 11994
rect 16689 11942 16719 11994
rect 16743 11942 16753 11994
rect 16753 11942 16799 11994
rect 16503 11940 16559 11942
rect 16583 11940 16639 11942
rect 16663 11940 16719 11942
rect 16743 11940 16799 11942
rect 14560 9274 14616 9276
rect 14640 9274 14696 9276
rect 14720 9274 14776 9276
rect 14800 9274 14856 9276
rect 14560 9222 14606 9274
rect 14606 9222 14616 9274
rect 14640 9222 14670 9274
rect 14670 9222 14682 9274
rect 14682 9222 14696 9274
rect 14720 9222 14734 9274
rect 14734 9222 14746 9274
rect 14746 9222 14776 9274
rect 14800 9222 14810 9274
rect 14810 9222 14856 9274
rect 14560 9220 14616 9222
rect 14640 9220 14696 9222
rect 14720 9220 14776 9222
rect 14800 9220 14856 9222
rect 14560 8186 14616 8188
rect 14640 8186 14696 8188
rect 14720 8186 14776 8188
rect 14800 8186 14856 8188
rect 14560 8134 14606 8186
rect 14606 8134 14616 8186
rect 14640 8134 14670 8186
rect 14670 8134 14682 8186
rect 14682 8134 14696 8186
rect 14720 8134 14734 8186
rect 14734 8134 14746 8186
rect 14746 8134 14776 8186
rect 14800 8134 14810 8186
rect 14810 8134 14856 8186
rect 14560 8132 14616 8134
rect 14640 8132 14696 8134
rect 14720 8132 14776 8134
rect 14800 8132 14856 8134
rect 14560 7098 14616 7100
rect 14640 7098 14696 7100
rect 14720 7098 14776 7100
rect 14800 7098 14856 7100
rect 14560 7046 14606 7098
rect 14606 7046 14616 7098
rect 14640 7046 14670 7098
rect 14670 7046 14682 7098
rect 14682 7046 14696 7098
rect 14720 7046 14734 7098
rect 14734 7046 14746 7098
rect 14746 7046 14776 7098
rect 14800 7046 14810 7098
rect 14810 7046 14856 7098
rect 14560 7044 14616 7046
rect 14640 7044 14696 7046
rect 14720 7044 14776 7046
rect 14800 7044 14856 7046
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 14560 6010 14616 6012
rect 14640 6010 14696 6012
rect 14720 6010 14776 6012
rect 14800 6010 14856 6012
rect 14560 5958 14606 6010
rect 14606 5958 14616 6010
rect 14640 5958 14670 6010
rect 14670 5958 14682 6010
rect 14682 5958 14696 6010
rect 14720 5958 14734 6010
rect 14734 5958 14746 6010
rect 14746 5958 14776 6010
rect 14800 5958 14810 6010
rect 14810 5958 14856 6010
rect 14560 5956 14616 5958
rect 14640 5956 14696 5958
rect 14720 5956 14776 5958
rect 14800 5956 14856 5958
rect 14560 4922 14616 4924
rect 14640 4922 14696 4924
rect 14720 4922 14776 4924
rect 14800 4922 14856 4924
rect 14560 4870 14606 4922
rect 14606 4870 14616 4922
rect 14640 4870 14670 4922
rect 14670 4870 14682 4922
rect 14682 4870 14696 4922
rect 14720 4870 14734 4922
rect 14734 4870 14746 4922
rect 14746 4870 14776 4922
rect 14800 4870 14810 4922
rect 14810 4870 14856 4922
rect 14560 4868 14616 4870
rect 14640 4868 14696 4870
rect 14720 4868 14776 4870
rect 14800 4868 14856 4870
rect 16503 10906 16559 10908
rect 16583 10906 16639 10908
rect 16663 10906 16719 10908
rect 16743 10906 16799 10908
rect 16503 10854 16549 10906
rect 16549 10854 16559 10906
rect 16583 10854 16613 10906
rect 16613 10854 16625 10906
rect 16625 10854 16639 10906
rect 16663 10854 16677 10906
rect 16677 10854 16689 10906
rect 16689 10854 16719 10906
rect 16743 10854 16753 10906
rect 16753 10854 16799 10906
rect 16503 10852 16559 10854
rect 16583 10852 16639 10854
rect 16663 10852 16719 10854
rect 16743 10852 16799 10854
rect 16503 9818 16559 9820
rect 16583 9818 16639 9820
rect 16663 9818 16719 9820
rect 16743 9818 16799 9820
rect 16503 9766 16549 9818
rect 16549 9766 16559 9818
rect 16583 9766 16613 9818
rect 16613 9766 16625 9818
rect 16625 9766 16639 9818
rect 16663 9766 16677 9818
rect 16677 9766 16689 9818
rect 16689 9766 16719 9818
rect 16743 9766 16753 9818
rect 16753 9766 16799 9818
rect 16503 9764 16559 9766
rect 16583 9764 16639 9766
rect 16663 9764 16719 9766
rect 16743 9764 16799 9766
rect 16302 9580 16358 9616
rect 16302 9560 16304 9580
rect 16304 9560 16356 9580
rect 16356 9560 16358 9580
rect 16503 8730 16559 8732
rect 16583 8730 16639 8732
rect 16663 8730 16719 8732
rect 16743 8730 16799 8732
rect 16503 8678 16549 8730
rect 16549 8678 16559 8730
rect 16583 8678 16613 8730
rect 16613 8678 16625 8730
rect 16625 8678 16639 8730
rect 16663 8678 16677 8730
rect 16677 8678 16689 8730
rect 16689 8678 16719 8730
rect 16743 8678 16753 8730
rect 16753 8678 16799 8730
rect 16503 8676 16559 8678
rect 16583 8676 16639 8678
rect 16663 8676 16719 8678
rect 16743 8676 16799 8678
rect 16503 7642 16559 7644
rect 16583 7642 16639 7644
rect 16663 7642 16719 7644
rect 16743 7642 16799 7644
rect 16503 7590 16549 7642
rect 16549 7590 16559 7642
rect 16583 7590 16613 7642
rect 16613 7590 16625 7642
rect 16625 7590 16639 7642
rect 16663 7590 16677 7642
rect 16677 7590 16689 7642
rect 16689 7590 16719 7642
rect 16743 7590 16753 7642
rect 16753 7590 16799 7642
rect 16503 7588 16559 7590
rect 16583 7588 16639 7590
rect 16663 7588 16719 7590
rect 16743 7588 16799 7590
rect 16503 6554 16559 6556
rect 16583 6554 16639 6556
rect 16663 6554 16719 6556
rect 16743 6554 16799 6556
rect 16503 6502 16549 6554
rect 16549 6502 16559 6554
rect 16583 6502 16613 6554
rect 16613 6502 16625 6554
rect 16625 6502 16639 6554
rect 16663 6502 16677 6554
rect 16677 6502 16689 6554
rect 16689 6502 16719 6554
rect 16743 6502 16753 6554
rect 16753 6502 16799 6554
rect 16503 6500 16559 6502
rect 16583 6500 16639 6502
rect 16663 6500 16719 6502
rect 16743 6500 16799 6502
rect 16946 5480 17002 5536
rect 16503 5466 16559 5468
rect 16583 5466 16639 5468
rect 16663 5466 16719 5468
rect 16743 5466 16799 5468
rect 16503 5414 16549 5466
rect 16549 5414 16559 5466
rect 16583 5414 16613 5466
rect 16613 5414 16625 5466
rect 16625 5414 16639 5466
rect 16663 5414 16677 5466
rect 16677 5414 16689 5466
rect 16689 5414 16719 5466
rect 16743 5414 16753 5466
rect 16753 5414 16799 5466
rect 16503 5412 16559 5414
rect 16583 5412 16639 5414
rect 16663 5412 16719 5414
rect 16743 5412 16799 5414
rect 16503 4378 16559 4380
rect 16583 4378 16639 4380
rect 16663 4378 16719 4380
rect 16743 4378 16799 4380
rect 16503 4326 16549 4378
rect 16549 4326 16559 4378
rect 16583 4326 16613 4378
rect 16613 4326 16625 4378
rect 16625 4326 16639 4378
rect 16663 4326 16677 4378
rect 16677 4326 16689 4378
rect 16689 4326 16719 4378
rect 16743 4326 16753 4378
rect 16753 4326 16799 4378
rect 16503 4324 16559 4326
rect 16583 4324 16639 4326
rect 16663 4324 16719 4326
rect 16743 4324 16799 4326
rect 14560 3834 14616 3836
rect 14640 3834 14696 3836
rect 14720 3834 14776 3836
rect 14800 3834 14856 3836
rect 14560 3782 14606 3834
rect 14606 3782 14616 3834
rect 14640 3782 14670 3834
rect 14670 3782 14682 3834
rect 14682 3782 14696 3834
rect 14720 3782 14734 3834
rect 14734 3782 14746 3834
rect 14746 3782 14776 3834
rect 14800 3782 14810 3834
rect 14810 3782 14856 3834
rect 14560 3780 14616 3782
rect 14640 3780 14696 3782
rect 14720 3780 14776 3782
rect 14800 3780 14856 3782
rect 14560 2746 14616 2748
rect 14640 2746 14696 2748
rect 14720 2746 14776 2748
rect 14800 2746 14856 2748
rect 14560 2694 14606 2746
rect 14606 2694 14616 2746
rect 14640 2694 14670 2746
rect 14670 2694 14682 2746
rect 14682 2694 14696 2746
rect 14720 2694 14734 2746
rect 14734 2694 14746 2746
rect 14746 2694 14776 2746
rect 14800 2694 14810 2746
rect 14810 2694 14856 2746
rect 14560 2692 14616 2694
rect 14640 2692 14696 2694
rect 14720 2692 14776 2694
rect 14800 2692 14856 2694
rect 16503 3290 16559 3292
rect 16583 3290 16639 3292
rect 16663 3290 16719 3292
rect 16743 3290 16799 3292
rect 16503 3238 16549 3290
rect 16549 3238 16559 3290
rect 16583 3238 16613 3290
rect 16613 3238 16625 3290
rect 16625 3238 16639 3290
rect 16663 3238 16677 3290
rect 16677 3238 16689 3290
rect 16689 3238 16719 3290
rect 16743 3238 16753 3290
rect 16753 3238 16799 3290
rect 16503 3236 16559 3238
rect 16583 3236 16639 3238
rect 16663 3236 16719 3238
rect 16743 3236 16799 3238
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 16503 2202 16559 2204
rect 16583 2202 16639 2204
rect 16663 2202 16719 2204
rect 16743 2202 16799 2204
rect 16503 2150 16549 2202
rect 16549 2150 16559 2202
rect 16583 2150 16613 2202
rect 16613 2150 16625 2202
rect 16625 2150 16639 2202
rect 16663 2150 16677 2202
rect 16677 2150 16689 2202
rect 16689 2150 16719 2202
rect 16743 2150 16753 2202
rect 16753 2150 16799 2202
rect 16503 2148 16559 2150
rect 16583 2148 16639 2150
rect 16663 2148 16719 2150
rect 16743 2148 16799 2150
rect 16486 1400 16542 1456
<< metal3 >>
rect 15929 17778 15995 17781
rect 17001 17778 17801 17808
rect 15929 17776 17801 17778
rect 15929 17720 15934 17776
rect 15990 17720 17801 17776
rect 15929 17718 17801 17720
rect 15929 17715 15995 17718
rect 17001 17688 17801 17718
rect 4832 17440 5148 17441
rect 4832 17376 4838 17440
rect 4902 17376 4918 17440
rect 4982 17376 4998 17440
rect 5062 17376 5078 17440
rect 5142 17376 5148 17440
rect 4832 17375 5148 17376
rect 8719 17440 9035 17441
rect 8719 17376 8725 17440
rect 8789 17376 8805 17440
rect 8869 17376 8885 17440
rect 8949 17376 8965 17440
rect 9029 17376 9035 17440
rect 8719 17375 9035 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 16493 17440 16809 17441
rect 16493 17376 16499 17440
rect 16563 17376 16579 17440
rect 16643 17376 16659 17440
rect 16723 17376 16739 17440
rect 16803 17376 16809 17440
rect 16493 17375 16809 17376
rect 2889 16896 3205 16897
rect 2889 16832 2895 16896
rect 2959 16832 2975 16896
rect 3039 16832 3055 16896
rect 3119 16832 3135 16896
rect 3199 16832 3205 16896
rect 2889 16831 3205 16832
rect 6776 16896 7092 16897
rect 6776 16832 6782 16896
rect 6846 16832 6862 16896
rect 6926 16832 6942 16896
rect 7006 16832 7022 16896
rect 7086 16832 7092 16896
rect 6776 16831 7092 16832
rect 10663 16896 10979 16897
rect 10663 16832 10669 16896
rect 10733 16832 10749 16896
rect 10813 16832 10829 16896
rect 10893 16832 10909 16896
rect 10973 16832 10979 16896
rect 10663 16831 10979 16832
rect 14550 16896 14866 16897
rect 14550 16832 14556 16896
rect 14620 16832 14636 16896
rect 14700 16832 14716 16896
rect 14780 16832 14796 16896
rect 14860 16832 14866 16896
rect 14550 16831 14866 16832
rect 0 16418 800 16448
rect 933 16418 999 16421
rect 0 16416 999 16418
rect 0 16360 938 16416
rect 994 16360 999 16416
rect 0 16358 999 16360
rect 0 16328 800 16358
rect 933 16355 999 16358
rect 4832 16352 5148 16353
rect 4832 16288 4838 16352
rect 4902 16288 4918 16352
rect 4982 16288 4998 16352
rect 5062 16288 5078 16352
rect 5142 16288 5148 16352
rect 4832 16287 5148 16288
rect 8719 16352 9035 16353
rect 8719 16288 8725 16352
rect 8789 16288 8805 16352
rect 8869 16288 8885 16352
rect 8949 16288 8965 16352
rect 9029 16288 9035 16352
rect 8719 16287 9035 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 16493 16352 16809 16353
rect 16493 16288 16499 16352
rect 16563 16288 16579 16352
rect 16643 16288 16659 16352
rect 16723 16288 16739 16352
rect 16803 16288 16809 16352
rect 16493 16287 16809 16288
rect 2889 15808 3205 15809
rect 2889 15744 2895 15808
rect 2959 15744 2975 15808
rect 3039 15744 3055 15808
rect 3119 15744 3135 15808
rect 3199 15744 3205 15808
rect 2889 15743 3205 15744
rect 6776 15808 7092 15809
rect 6776 15744 6782 15808
rect 6846 15744 6862 15808
rect 6926 15744 6942 15808
rect 7006 15744 7022 15808
rect 7086 15744 7092 15808
rect 6776 15743 7092 15744
rect 10663 15808 10979 15809
rect 10663 15744 10669 15808
rect 10733 15744 10749 15808
rect 10813 15744 10829 15808
rect 10893 15744 10909 15808
rect 10973 15744 10979 15808
rect 10663 15743 10979 15744
rect 14550 15808 14866 15809
rect 14550 15744 14556 15808
rect 14620 15744 14636 15808
rect 14700 15744 14716 15808
rect 14780 15744 14796 15808
rect 14860 15744 14866 15808
rect 14550 15743 14866 15744
rect 4832 15264 5148 15265
rect 4832 15200 4838 15264
rect 4902 15200 4918 15264
rect 4982 15200 4998 15264
rect 5062 15200 5078 15264
rect 5142 15200 5148 15264
rect 4832 15199 5148 15200
rect 8719 15264 9035 15265
rect 8719 15200 8725 15264
rect 8789 15200 8805 15264
rect 8869 15200 8885 15264
rect 8949 15200 8965 15264
rect 9029 15200 9035 15264
rect 8719 15199 9035 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 16493 15264 16809 15265
rect 16493 15200 16499 15264
rect 16563 15200 16579 15264
rect 16643 15200 16659 15264
rect 16723 15200 16739 15264
rect 16803 15200 16809 15264
rect 16493 15199 16809 15200
rect 2889 14720 3205 14721
rect 2889 14656 2895 14720
rect 2959 14656 2975 14720
rect 3039 14656 3055 14720
rect 3119 14656 3135 14720
rect 3199 14656 3205 14720
rect 2889 14655 3205 14656
rect 6776 14720 7092 14721
rect 6776 14656 6782 14720
rect 6846 14656 6862 14720
rect 6926 14656 6942 14720
rect 7006 14656 7022 14720
rect 7086 14656 7092 14720
rect 6776 14655 7092 14656
rect 10663 14720 10979 14721
rect 10663 14656 10669 14720
rect 10733 14656 10749 14720
rect 10813 14656 10829 14720
rect 10893 14656 10909 14720
rect 10973 14656 10979 14720
rect 10663 14655 10979 14656
rect 14550 14720 14866 14721
rect 14550 14656 14556 14720
rect 14620 14656 14636 14720
rect 14700 14656 14716 14720
rect 14780 14656 14796 14720
rect 14860 14656 14866 14720
rect 14550 14655 14866 14656
rect 4832 14176 5148 14177
rect 4832 14112 4838 14176
rect 4902 14112 4918 14176
rect 4982 14112 4998 14176
rect 5062 14112 5078 14176
rect 5142 14112 5148 14176
rect 4832 14111 5148 14112
rect 8719 14176 9035 14177
rect 8719 14112 8725 14176
rect 8789 14112 8805 14176
rect 8869 14112 8885 14176
rect 8949 14112 8965 14176
rect 9029 14112 9035 14176
rect 8719 14111 9035 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 16493 14176 16809 14177
rect 16493 14112 16499 14176
rect 16563 14112 16579 14176
rect 16643 14112 16659 14176
rect 16723 14112 16739 14176
rect 16803 14112 16809 14176
rect 16493 14111 16809 14112
rect 16573 13698 16639 13701
rect 17001 13698 17801 13728
rect 16573 13696 17801 13698
rect 16573 13640 16578 13696
rect 16634 13640 17801 13696
rect 16573 13638 17801 13640
rect 16573 13635 16639 13638
rect 2889 13632 3205 13633
rect 2889 13568 2895 13632
rect 2959 13568 2975 13632
rect 3039 13568 3055 13632
rect 3119 13568 3135 13632
rect 3199 13568 3205 13632
rect 2889 13567 3205 13568
rect 6776 13632 7092 13633
rect 6776 13568 6782 13632
rect 6846 13568 6862 13632
rect 6926 13568 6942 13632
rect 7006 13568 7022 13632
rect 7086 13568 7092 13632
rect 6776 13567 7092 13568
rect 10663 13632 10979 13633
rect 10663 13568 10669 13632
rect 10733 13568 10749 13632
rect 10813 13568 10829 13632
rect 10893 13568 10909 13632
rect 10973 13568 10979 13632
rect 10663 13567 10979 13568
rect 14550 13632 14866 13633
rect 14550 13568 14556 13632
rect 14620 13568 14636 13632
rect 14700 13568 14716 13632
rect 14780 13568 14796 13632
rect 14860 13568 14866 13632
rect 17001 13608 17801 13638
rect 14550 13567 14866 13568
rect 4832 13088 5148 13089
rect 4832 13024 4838 13088
rect 4902 13024 4918 13088
rect 4982 13024 4998 13088
rect 5062 13024 5078 13088
rect 5142 13024 5148 13088
rect 4832 13023 5148 13024
rect 8719 13088 9035 13089
rect 8719 13024 8725 13088
rect 8789 13024 8805 13088
rect 8869 13024 8885 13088
rect 8949 13024 8965 13088
rect 9029 13024 9035 13088
rect 8719 13023 9035 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 16493 13088 16809 13089
rect 16493 13024 16499 13088
rect 16563 13024 16579 13088
rect 16643 13024 16659 13088
rect 16723 13024 16739 13088
rect 16803 13024 16809 13088
rect 16493 13023 16809 13024
rect 5441 12746 5507 12749
rect 9857 12746 9923 12749
rect 5441 12744 9923 12746
rect 5441 12688 5446 12744
rect 5502 12688 9862 12744
rect 9918 12688 9923 12744
rect 5441 12686 9923 12688
rect 5441 12683 5507 12686
rect 9857 12683 9923 12686
rect 2889 12544 3205 12545
rect 2889 12480 2895 12544
rect 2959 12480 2975 12544
rect 3039 12480 3055 12544
rect 3119 12480 3135 12544
rect 3199 12480 3205 12544
rect 2889 12479 3205 12480
rect 6776 12544 7092 12545
rect 6776 12480 6782 12544
rect 6846 12480 6862 12544
rect 6926 12480 6942 12544
rect 7006 12480 7022 12544
rect 7086 12480 7092 12544
rect 6776 12479 7092 12480
rect 10663 12544 10979 12545
rect 10663 12480 10669 12544
rect 10733 12480 10749 12544
rect 10813 12480 10829 12544
rect 10893 12480 10909 12544
rect 10973 12480 10979 12544
rect 10663 12479 10979 12480
rect 14550 12544 14866 12545
rect 14550 12480 14556 12544
rect 14620 12480 14636 12544
rect 14700 12480 14716 12544
rect 14780 12480 14796 12544
rect 14860 12480 14866 12544
rect 14550 12479 14866 12480
rect 0 12338 800 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 4832 12000 5148 12001
rect 4832 11936 4838 12000
rect 4902 11936 4918 12000
rect 4982 11936 4998 12000
rect 5062 11936 5078 12000
rect 5142 11936 5148 12000
rect 4832 11935 5148 11936
rect 8719 12000 9035 12001
rect 8719 11936 8725 12000
rect 8789 11936 8805 12000
rect 8869 11936 8885 12000
rect 8949 11936 8965 12000
rect 9029 11936 9035 12000
rect 8719 11935 9035 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 16493 12000 16809 12001
rect 16493 11936 16499 12000
rect 16563 11936 16579 12000
rect 16643 11936 16659 12000
rect 16723 11936 16739 12000
rect 16803 11936 16809 12000
rect 16493 11935 16809 11936
rect 2889 11456 3205 11457
rect 2889 11392 2895 11456
rect 2959 11392 2975 11456
rect 3039 11392 3055 11456
rect 3119 11392 3135 11456
rect 3199 11392 3205 11456
rect 2889 11391 3205 11392
rect 6776 11456 7092 11457
rect 6776 11392 6782 11456
rect 6846 11392 6862 11456
rect 6926 11392 6942 11456
rect 7006 11392 7022 11456
rect 7086 11392 7092 11456
rect 6776 11391 7092 11392
rect 10663 11456 10979 11457
rect 10663 11392 10669 11456
rect 10733 11392 10749 11456
rect 10813 11392 10829 11456
rect 10893 11392 10909 11456
rect 10973 11392 10979 11456
rect 10663 11391 10979 11392
rect 14550 11456 14866 11457
rect 14550 11392 14556 11456
rect 14620 11392 14636 11456
rect 14700 11392 14716 11456
rect 14780 11392 14796 11456
rect 14860 11392 14866 11456
rect 14550 11391 14866 11392
rect 4832 10912 5148 10913
rect 4832 10848 4838 10912
rect 4902 10848 4918 10912
rect 4982 10848 4998 10912
rect 5062 10848 5078 10912
rect 5142 10848 5148 10912
rect 4832 10847 5148 10848
rect 8719 10912 9035 10913
rect 8719 10848 8725 10912
rect 8789 10848 8805 10912
rect 8869 10848 8885 10912
rect 8949 10848 8965 10912
rect 9029 10848 9035 10912
rect 8719 10847 9035 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 16493 10912 16809 10913
rect 16493 10848 16499 10912
rect 16563 10848 16579 10912
rect 16643 10848 16659 10912
rect 16723 10848 16739 10912
rect 16803 10848 16809 10912
rect 16493 10847 16809 10848
rect 2889 10368 3205 10369
rect 2889 10304 2895 10368
rect 2959 10304 2975 10368
rect 3039 10304 3055 10368
rect 3119 10304 3135 10368
rect 3199 10304 3205 10368
rect 2889 10303 3205 10304
rect 6776 10368 7092 10369
rect 6776 10304 6782 10368
rect 6846 10304 6862 10368
rect 6926 10304 6942 10368
rect 7006 10304 7022 10368
rect 7086 10304 7092 10368
rect 6776 10303 7092 10304
rect 10663 10368 10979 10369
rect 10663 10304 10669 10368
rect 10733 10304 10749 10368
rect 10813 10304 10829 10368
rect 10893 10304 10909 10368
rect 10973 10304 10979 10368
rect 10663 10303 10979 10304
rect 14550 10368 14866 10369
rect 14550 10304 14556 10368
rect 14620 10304 14636 10368
rect 14700 10304 14716 10368
rect 14780 10304 14796 10368
rect 14860 10304 14866 10368
rect 14550 10303 14866 10304
rect 4832 9824 5148 9825
rect 4832 9760 4838 9824
rect 4902 9760 4918 9824
rect 4982 9760 4998 9824
rect 5062 9760 5078 9824
rect 5142 9760 5148 9824
rect 4832 9759 5148 9760
rect 8719 9824 9035 9825
rect 8719 9760 8725 9824
rect 8789 9760 8805 9824
rect 8869 9760 8885 9824
rect 8949 9760 8965 9824
rect 9029 9760 9035 9824
rect 8719 9759 9035 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 16493 9824 16809 9825
rect 16493 9760 16499 9824
rect 16563 9760 16579 9824
rect 16643 9760 16659 9824
rect 16723 9760 16739 9824
rect 16803 9760 16809 9824
rect 16493 9759 16809 9760
rect 16297 9618 16363 9621
rect 17001 9618 17801 9648
rect 16297 9616 17801 9618
rect 16297 9560 16302 9616
rect 16358 9560 17801 9616
rect 16297 9558 17801 9560
rect 16297 9555 16363 9558
rect 17001 9528 17801 9558
rect 2889 9280 3205 9281
rect 2889 9216 2895 9280
rect 2959 9216 2975 9280
rect 3039 9216 3055 9280
rect 3119 9216 3135 9280
rect 3199 9216 3205 9280
rect 2889 9215 3205 9216
rect 6776 9280 7092 9281
rect 6776 9216 6782 9280
rect 6846 9216 6862 9280
rect 6926 9216 6942 9280
rect 7006 9216 7022 9280
rect 7086 9216 7092 9280
rect 6776 9215 7092 9216
rect 10663 9280 10979 9281
rect 10663 9216 10669 9280
rect 10733 9216 10749 9280
rect 10813 9216 10829 9280
rect 10893 9216 10909 9280
rect 10973 9216 10979 9280
rect 10663 9215 10979 9216
rect 14550 9280 14866 9281
rect 14550 9216 14556 9280
rect 14620 9216 14636 9280
rect 14700 9216 14716 9280
rect 14780 9216 14796 9280
rect 14860 9216 14866 9280
rect 14550 9215 14866 9216
rect 4832 8736 5148 8737
rect 4832 8672 4838 8736
rect 4902 8672 4918 8736
rect 4982 8672 4998 8736
rect 5062 8672 5078 8736
rect 5142 8672 5148 8736
rect 4832 8671 5148 8672
rect 8719 8736 9035 8737
rect 8719 8672 8725 8736
rect 8789 8672 8805 8736
rect 8869 8672 8885 8736
rect 8949 8672 8965 8736
rect 9029 8672 9035 8736
rect 8719 8671 9035 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 16493 8736 16809 8737
rect 16493 8672 16499 8736
rect 16563 8672 16579 8736
rect 16643 8672 16659 8736
rect 16723 8672 16739 8736
rect 16803 8672 16809 8736
rect 16493 8671 16809 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 2889 8192 3205 8193
rect 2889 8128 2895 8192
rect 2959 8128 2975 8192
rect 3039 8128 3055 8192
rect 3119 8128 3135 8192
rect 3199 8128 3205 8192
rect 2889 8127 3205 8128
rect 6776 8192 7092 8193
rect 6776 8128 6782 8192
rect 6846 8128 6862 8192
rect 6926 8128 6942 8192
rect 7006 8128 7022 8192
rect 7086 8128 7092 8192
rect 6776 8127 7092 8128
rect 10663 8192 10979 8193
rect 10663 8128 10669 8192
rect 10733 8128 10749 8192
rect 10813 8128 10829 8192
rect 10893 8128 10909 8192
rect 10973 8128 10979 8192
rect 10663 8127 10979 8128
rect 14550 8192 14866 8193
rect 14550 8128 14556 8192
rect 14620 8128 14636 8192
rect 14700 8128 14716 8192
rect 14780 8128 14796 8192
rect 14860 8128 14866 8192
rect 14550 8127 14866 8128
rect 4832 7648 5148 7649
rect 4832 7584 4838 7648
rect 4902 7584 4918 7648
rect 4982 7584 4998 7648
rect 5062 7584 5078 7648
rect 5142 7584 5148 7648
rect 4832 7583 5148 7584
rect 8719 7648 9035 7649
rect 8719 7584 8725 7648
rect 8789 7584 8805 7648
rect 8869 7584 8885 7648
rect 8949 7584 8965 7648
rect 9029 7584 9035 7648
rect 8719 7583 9035 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 16493 7648 16809 7649
rect 16493 7584 16499 7648
rect 16563 7584 16579 7648
rect 16643 7584 16659 7648
rect 16723 7584 16739 7648
rect 16803 7584 16809 7648
rect 16493 7583 16809 7584
rect 2889 7104 3205 7105
rect 2889 7040 2895 7104
rect 2959 7040 2975 7104
rect 3039 7040 3055 7104
rect 3119 7040 3135 7104
rect 3199 7040 3205 7104
rect 2889 7039 3205 7040
rect 6776 7104 7092 7105
rect 6776 7040 6782 7104
rect 6846 7040 6862 7104
rect 6926 7040 6942 7104
rect 7006 7040 7022 7104
rect 7086 7040 7092 7104
rect 6776 7039 7092 7040
rect 10663 7104 10979 7105
rect 10663 7040 10669 7104
rect 10733 7040 10749 7104
rect 10813 7040 10829 7104
rect 10893 7040 10909 7104
rect 10973 7040 10979 7104
rect 10663 7039 10979 7040
rect 14550 7104 14866 7105
rect 14550 7040 14556 7104
rect 14620 7040 14636 7104
rect 14700 7040 14716 7104
rect 14780 7040 14796 7104
rect 14860 7040 14866 7104
rect 14550 7039 14866 7040
rect 4832 6560 5148 6561
rect 4832 6496 4838 6560
rect 4902 6496 4918 6560
rect 4982 6496 4998 6560
rect 5062 6496 5078 6560
rect 5142 6496 5148 6560
rect 4832 6495 5148 6496
rect 8719 6560 9035 6561
rect 8719 6496 8725 6560
rect 8789 6496 8805 6560
rect 8869 6496 8885 6560
rect 8949 6496 8965 6560
rect 9029 6496 9035 6560
rect 8719 6495 9035 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 16493 6560 16809 6561
rect 16493 6496 16499 6560
rect 16563 6496 16579 6560
rect 16643 6496 16659 6560
rect 16723 6496 16739 6560
rect 16803 6496 16809 6560
rect 16493 6495 16809 6496
rect 2889 6016 3205 6017
rect 2889 5952 2895 6016
rect 2959 5952 2975 6016
rect 3039 5952 3055 6016
rect 3119 5952 3135 6016
rect 3199 5952 3205 6016
rect 2889 5951 3205 5952
rect 6776 6016 7092 6017
rect 6776 5952 6782 6016
rect 6846 5952 6862 6016
rect 6926 5952 6942 6016
rect 7006 5952 7022 6016
rect 7086 5952 7092 6016
rect 6776 5951 7092 5952
rect 10663 6016 10979 6017
rect 10663 5952 10669 6016
rect 10733 5952 10749 6016
rect 10813 5952 10829 6016
rect 10893 5952 10909 6016
rect 10973 5952 10979 6016
rect 10663 5951 10979 5952
rect 14550 6016 14866 6017
rect 14550 5952 14556 6016
rect 14620 5952 14636 6016
rect 14700 5952 14716 6016
rect 14780 5952 14796 6016
rect 14860 5952 14866 6016
rect 14550 5951 14866 5952
rect 17001 5541 17801 5568
rect 16941 5536 17801 5541
rect 16941 5480 16946 5536
rect 17002 5480 17801 5536
rect 16941 5475 17801 5480
rect 4832 5472 5148 5473
rect 4832 5408 4838 5472
rect 4902 5408 4918 5472
rect 4982 5408 4998 5472
rect 5062 5408 5078 5472
rect 5142 5408 5148 5472
rect 4832 5407 5148 5408
rect 8719 5472 9035 5473
rect 8719 5408 8725 5472
rect 8789 5408 8805 5472
rect 8869 5408 8885 5472
rect 8949 5408 8965 5472
rect 9029 5408 9035 5472
rect 8719 5407 9035 5408
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 16493 5472 16809 5473
rect 16493 5408 16499 5472
rect 16563 5408 16579 5472
rect 16643 5408 16659 5472
rect 16723 5408 16739 5472
rect 16803 5408 16809 5472
rect 17001 5448 17801 5475
rect 16493 5407 16809 5408
rect 2889 4928 3205 4929
rect 2889 4864 2895 4928
rect 2959 4864 2975 4928
rect 3039 4864 3055 4928
rect 3119 4864 3135 4928
rect 3199 4864 3205 4928
rect 2889 4863 3205 4864
rect 6776 4928 7092 4929
rect 6776 4864 6782 4928
rect 6846 4864 6862 4928
rect 6926 4864 6942 4928
rect 7006 4864 7022 4928
rect 7086 4864 7092 4928
rect 6776 4863 7092 4864
rect 10663 4928 10979 4929
rect 10663 4864 10669 4928
rect 10733 4864 10749 4928
rect 10813 4864 10829 4928
rect 10893 4864 10909 4928
rect 10973 4864 10979 4928
rect 10663 4863 10979 4864
rect 14550 4928 14866 4929
rect 14550 4864 14556 4928
rect 14620 4864 14636 4928
rect 14700 4864 14716 4928
rect 14780 4864 14796 4928
rect 14860 4864 14866 4928
rect 14550 4863 14866 4864
rect 4832 4384 5148 4385
rect 4832 4320 4838 4384
rect 4902 4320 4918 4384
rect 4982 4320 4998 4384
rect 5062 4320 5078 4384
rect 5142 4320 5148 4384
rect 4832 4319 5148 4320
rect 8719 4384 9035 4385
rect 8719 4320 8725 4384
rect 8789 4320 8805 4384
rect 8869 4320 8885 4384
rect 8949 4320 8965 4384
rect 9029 4320 9035 4384
rect 8719 4319 9035 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 16493 4384 16809 4385
rect 16493 4320 16499 4384
rect 16563 4320 16579 4384
rect 16643 4320 16659 4384
rect 16723 4320 16739 4384
rect 16803 4320 16809 4384
rect 16493 4319 16809 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 2889 3840 3205 3841
rect 2889 3776 2895 3840
rect 2959 3776 2975 3840
rect 3039 3776 3055 3840
rect 3119 3776 3135 3840
rect 3199 3776 3205 3840
rect 2889 3775 3205 3776
rect 6776 3840 7092 3841
rect 6776 3776 6782 3840
rect 6846 3776 6862 3840
rect 6926 3776 6942 3840
rect 7006 3776 7022 3840
rect 7086 3776 7092 3840
rect 6776 3775 7092 3776
rect 10663 3840 10979 3841
rect 10663 3776 10669 3840
rect 10733 3776 10749 3840
rect 10813 3776 10829 3840
rect 10893 3776 10909 3840
rect 10973 3776 10979 3840
rect 10663 3775 10979 3776
rect 14550 3840 14866 3841
rect 14550 3776 14556 3840
rect 14620 3776 14636 3840
rect 14700 3776 14716 3840
rect 14780 3776 14796 3840
rect 14860 3776 14866 3840
rect 14550 3775 14866 3776
rect 4832 3296 5148 3297
rect 4832 3232 4838 3296
rect 4902 3232 4918 3296
rect 4982 3232 4998 3296
rect 5062 3232 5078 3296
rect 5142 3232 5148 3296
rect 4832 3231 5148 3232
rect 8719 3296 9035 3297
rect 8719 3232 8725 3296
rect 8789 3232 8805 3296
rect 8869 3232 8885 3296
rect 8949 3232 8965 3296
rect 9029 3232 9035 3296
rect 8719 3231 9035 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 16493 3296 16809 3297
rect 16493 3232 16499 3296
rect 16563 3232 16579 3296
rect 16643 3232 16659 3296
rect 16723 3232 16739 3296
rect 16803 3232 16809 3296
rect 16493 3231 16809 3232
rect 2889 2752 3205 2753
rect 2889 2688 2895 2752
rect 2959 2688 2975 2752
rect 3039 2688 3055 2752
rect 3119 2688 3135 2752
rect 3199 2688 3205 2752
rect 2889 2687 3205 2688
rect 6776 2752 7092 2753
rect 6776 2688 6782 2752
rect 6846 2688 6862 2752
rect 6926 2688 6942 2752
rect 7006 2688 7022 2752
rect 7086 2688 7092 2752
rect 6776 2687 7092 2688
rect 10663 2752 10979 2753
rect 10663 2688 10669 2752
rect 10733 2688 10749 2752
rect 10813 2688 10829 2752
rect 10893 2688 10909 2752
rect 10973 2688 10979 2752
rect 10663 2687 10979 2688
rect 14550 2752 14866 2753
rect 14550 2688 14556 2752
rect 14620 2688 14636 2752
rect 14700 2688 14716 2752
rect 14780 2688 14796 2752
rect 14860 2688 14866 2752
rect 14550 2687 14866 2688
rect 4832 2208 5148 2209
rect 4832 2144 4838 2208
rect 4902 2144 4918 2208
rect 4982 2144 4998 2208
rect 5062 2144 5078 2208
rect 5142 2144 5148 2208
rect 4832 2143 5148 2144
rect 8719 2208 9035 2209
rect 8719 2144 8725 2208
rect 8789 2144 8805 2208
rect 8869 2144 8885 2208
rect 8949 2144 8965 2208
rect 9029 2144 9035 2208
rect 8719 2143 9035 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 16493 2208 16809 2209
rect 16493 2144 16499 2208
rect 16563 2144 16579 2208
rect 16643 2144 16659 2208
rect 16723 2144 16739 2208
rect 16803 2144 16809 2208
rect 16493 2143 16809 2144
rect 16481 1458 16547 1461
rect 17001 1458 17801 1488
rect 16481 1456 17801 1458
rect 16481 1400 16486 1456
rect 16542 1400 17801 1456
rect 16481 1398 17801 1400
rect 16481 1395 16547 1398
rect 17001 1368 17801 1398
<< via3 >>
rect 4838 17436 4902 17440
rect 4838 17380 4842 17436
rect 4842 17380 4898 17436
rect 4898 17380 4902 17436
rect 4838 17376 4902 17380
rect 4918 17436 4982 17440
rect 4918 17380 4922 17436
rect 4922 17380 4978 17436
rect 4978 17380 4982 17436
rect 4918 17376 4982 17380
rect 4998 17436 5062 17440
rect 4998 17380 5002 17436
rect 5002 17380 5058 17436
rect 5058 17380 5062 17436
rect 4998 17376 5062 17380
rect 5078 17436 5142 17440
rect 5078 17380 5082 17436
rect 5082 17380 5138 17436
rect 5138 17380 5142 17436
rect 5078 17376 5142 17380
rect 8725 17436 8789 17440
rect 8725 17380 8729 17436
rect 8729 17380 8785 17436
rect 8785 17380 8789 17436
rect 8725 17376 8789 17380
rect 8805 17436 8869 17440
rect 8805 17380 8809 17436
rect 8809 17380 8865 17436
rect 8865 17380 8869 17436
rect 8805 17376 8869 17380
rect 8885 17436 8949 17440
rect 8885 17380 8889 17436
rect 8889 17380 8945 17436
rect 8945 17380 8949 17436
rect 8885 17376 8949 17380
rect 8965 17436 9029 17440
rect 8965 17380 8969 17436
rect 8969 17380 9025 17436
rect 9025 17380 9029 17436
rect 8965 17376 9029 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 16499 17436 16563 17440
rect 16499 17380 16503 17436
rect 16503 17380 16559 17436
rect 16559 17380 16563 17436
rect 16499 17376 16563 17380
rect 16579 17436 16643 17440
rect 16579 17380 16583 17436
rect 16583 17380 16639 17436
rect 16639 17380 16643 17436
rect 16579 17376 16643 17380
rect 16659 17436 16723 17440
rect 16659 17380 16663 17436
rect 16663 17380 16719 17436
rect 16719 17380 16723 17436
rect 16659 17376 16723 17380
rect 16739 17436 16803 17440
rect 16739 17380 16743 17436
rect 16743 17380 16799 17436
rect 16799 17380 16803 17436
rect 16739 17376 16803 17380
rect 2895 16892 2959 16896
rect 2895 16836 2899 16892
rect 2899 16836 2955 16892
rect 2955 16836 2959 16892
rect 2895 16832 2959 16836
rect 2975 16892 3039 16896
rect 2975 16836 2979 16892
rect 2979 16836 3035 16892
rect 3035 16836 3039 16892
rect 2975 16832 3039 16836
rect 3055 16892 3119 16896
rect 3055 16836 3059 16892
rect 3059 16836 3115 16892
rect 3115 16836 3119 16892
rect 3055 16832 3119 16836
rect 3135 16892 3199 16896
rect 3135 16836 3139 16892
rect 3139 16836 3195 16892
rect 3195 16836 3199 16892
rect 3135 16832 3199 16836
rect 6782 16892 6846 16896
rect 6782 16836 6786 16892
rect 6786 16836 6842 16892
rect 6842 16836 6846 16892
rect 6782 16832 6846 16836
rect 6862 16892 6926 16896
rect 6862 16836 6866 16892
rect 6866 16836 6922 16892
rect 6922 16836 6926 16892
rect 6862 16832 6926 16836
rect 6942 16892 7006 16896
rect 6942 16836 6946 16892
rect 6946 16836 7002 16892
rect 7002 16836 7006 16892
rect 6942 16832 7006 16836
rect 7022 16892 7086 16896
rect 7022 16836 7026 16892
rect 7026 16836 7082 16892
rect 7082 16836 7086 16892
rect 7022 16832 7086 16836
rect 10669 16892 10733 16896
rect 10669 16836 10673 16892
rect 10673 16836 10729 16892
rect 10729 16836 10733 16892
rect 10669 16832 10733 16836
rect 10749 16892 10813 16896
rect 10749 16836 10753 16892
rect 10753 16836 10809 16892
rect 10809 16836 10813 16892
rect 10749 16832 10813 16836
rect 10829 16892 10893 16896
rect 10829 16836 10833 16892
rect 10833 16836 10889 16892
rect 10889 16836 10893 16892
rect 10829 16832 10893 16836
rect 10909 16892 10973 16896
rect 10909 16836 10913 16892
rect 10913 16836 10969 16892
rect 10969 16836 10973 16892
rect 10909 16832 10973 16836
rect 14556 16892 14620 16896
rect 14556 16836 14560 16892
rect 14560 16836 14616 16892
rect 14616 16836 14620 16892
rect 14556 16832 14620 16836
rect 14636 16892 14700 16896
rect 14636 16836 14640 16892
rect 14640 16836 14696 16892
rect 14696 16836 14700 16892
rect 14636 16832 14700 16836
rect 14716 16892 14780 16896
rect 14716 16836 14720 16892
rect 14720 16836 14776 16892
rect 14776 16836 14780 16892
rect 14716 16832 14780 16836
rect 14796 16892 14860 16896
rect 14796 16836 14800 16892
rect 14800 16836 14856 16892
rect 14856 16836 14860 16892
rect 14796 16832 14860 16836
rect 4838 16348 4902 16352
rect 4838 16292 4842 16348
rect 4842 16292 4898 16348
rect 4898 16292 4902 16348
rect 4838 16288 4902 16292
rect 4918 16348 4982 16352
rect 4918 16292 4922 16348
rect 4922 16292 4978 16348
rect 4978 16292 4982 16348
rect 4918 16288 4982 16292
rect 4998 16348 5062 16352
rect 4998 16292 5002 16348
rect 5002 16292 5058 16348
rect 5058 16292 5062 16348
rect 4998 16288 5062 16292
rect 5078 16348 5142 16352
rect 5078 16292 5082 16348
rect 5082 16292 5138 16348
rect 5138 16292 5142 16348
rect 5078 16288 5142 16292
rect 8725 16348 8789 16352
rect 8725 16292 8729 16348
rect 8729 16292 8785 16348
rect 8785 16292 8789 16348
rect 8725 16288 8789 16292
rect 8805 16348 8869 16352
rect 8805 16292 8809 16348
rect 8809 16292 8865 16348
rect 8865 16292 8869 16348
rect 8805 16288 8869 16292
rect 8885 16348 8949 16352
rect 8885 16292 8889 16348
rect 8889 16292 8945 16348
rect 8945 16292 8949 16348
rect 8885 16288 8949 16292
rect 8965 16348 9029 16352
rect 8965 16292 8969 16348
rect 8969 16292 9025 16348
rect 9025 16292 9029 16348
rect 8965 16288 9029 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 16499 16348 16563 16352
rect 16499 16292 16503 16348
rect 16503 16292 16559 16348
rect 16559 16292 16563 16348
rect 16499 16288 16563 16292
rect 16579 16348 16643 16352
rect 16579 16292 16583 16348
rect 16583 16292 16639 16348
rect 16639 16292 16643 16348
rect 16579 16288 16643 16292
rect 16659 16348 16723 16352
rect 16659 16292 16663 16348
rect 16663 16292 16719 16348
rect 16719 16292 16723 16348
rect 16659 16288 16723 16292
rect 16739 16348 16803 16352
rect 16739 16292 16743 16348
rect 16743 16292 16799 16348
rect 16799 16292 16803 16348
rect 16739 16288 16803 16292
rect 2895 15804 2959 15808
rect 2895 15748 2899 15804
rect 2899 15748 2955 15804
rect 2955 15748 2959 15804
rect 2895 15744 2959 15748
rect 2975 15804 3039 15808
rect 2975 15748 2979 15804
rect 2979 15748 3035 15804
rect 3035 15748 3039 15804
rect 2975 15744 3039 15748
rect 3055 15804 3119 15808
rect 3055 15748 3059 15804
rect 3059 15748 3115 15804
rect 3115 15748 3119 15804
rect 3055 15744 3119 15748
rect 3135 15804 3199 15808
rect 3135 15748 3139 15804
rect 3139 15748 3195 15804
rect 3195 15748 3199 15804
rect 3135 15744 3199 15748
rect 6782 15804 6846 15808
rect 6782 15748 6786 15804
rect 6786 15748 6842 15804
rect 6842 15748 6846 15804
rect 6782 15744 6846 15748
rect 6862 15804 6926 15808
rect 6862 15748 6866 15804
rect 6866 15748 6922 15804
rect 6922 15748 6926 15804
rect 6862 15744 6926 15748
rect 6942 15804 7006 15808
rect 6942 15748 6946 15804
rect 6946 15748 7002 15804
rect 7002 15748 7006 15804
rect 6942 15744 7006 15748
rect 7022 15804 7086 15808
rect 7022 15748 7026 15804
rect 7026 15748 7082 15804
rect 7082 15748 7086 15804
rect 7022 15744 7086 15748
rect 10669 15804 10733 15808
rect 10669 15748 10673 15804
rect 10673 15748 10729 15804
rect 10729 15748 10733 15804
rect 10669 15744 10733 15748
rect 10749 15804 10813 15808
rect 10749 15748 10753 15804
rect 10753 15748 10809 15804
rect 10809 15748 10813 15804
rect 10749 15744 10813 15748
rect 10829 15804 10893 15808
rect 10829 15748 10833 15804
rect 10833 15748 10889 15804
rect 10889 15748 10893 15804
rect 10829 15744 10893 15748
rect 10909 15804 10973 15808
rect 10909 15748 10913 15804
rect 10913 15748 10969 15804
rect 10969 15748 10973 15804
rect 10909 15744 10973 15748
rect 14556 15804 14620 15808
rect 14556 15748 14560 15804
rect 14560 15748 14616 15804
rect 14616 15748 14620 15804
rect 14556 15744 14620 15748
rect 14636 15804 14700 15808
rect 14636 15748 14640 15804
rect 14640 15748 14696 15804
rect 14696 15748 14700 15804
rect 14636 15744 14700 15748
rect 14716 15804 14780 15808
rect 14716 15748 14720 15804
rect 14720 15748 14776 15804
rect 14776 15748 14780 15804
rect 14716 15744 14780 15748
rect 14796 15804 14860 15808
rect 14796 15748 14800 15804
rect 14800 15748 14856 15804
rect 14856 15748 14860 15804
rect 14796 15744 14860 15748
rect 4838 15260 4902 15264
rect 4838 15204 4842 15260
rect 4842 15204 4898 15260
rect 4898 15204 4902 15260
rect 4838 15200 4902 15204
rect 4918 15260 4982 15264
rect 4918 15204 4922 15260
rect 4922 15204 4978 15260
rect 4978 15204 4982 15260
rect 4918 15200 4982 15204
rect 4998 15260 5062 15264
rect 4998 15204 5002 15260
rect 5002 15204 5058 15260
rect 5058 15204 5062 15260
rect 4998 15200 5062 15204
rect 5078 15260 5142 15264
rect 5078 15204 5082 15260
rect 5082 15204 5138 15260
rect 5138 15204 5142 15260
rect 5078 15200 5142 15204
rect 8725 15260 8789 15264
rect 8725 15204 8729 15260
rect 8729 15204 8785 15260
rect 8785 15204 8789 15260
rect 8725 15200 8789 15204
rect 8805 15260 8869 15264
rect 8805 15204 8809 15260
rect 8809 15204 8865 15260
rect 8865 15204 8869 15260
rect 8805 15200 8869 15204
rect 8885 15260 8949 15264
rect 8885 15204 8889 15260
rect 8889 15204 8945 15260
rect 8945 15204 8949 15260
rect 8885 15200 8949 15204
rect 8965 15260 9029 15264
rect 8965 15204 8969 15260
rect 8969 15204 9025 15260
rect 9025 15204 9029 15260
rect 8965 15200 9029 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 16499 15260 16563 15264
rect 16499 15204 16503 15260
rect 16503 15204 16559 15260
rect 16559 15204 16563 15260
rect 16499 15200 16563 15204
rect 16579 15260 16643 15264
rect 16579 15204 16583 15260
rect 16583 15204 16639 15260
rect 16639 15204 16643 15260
rect 16579 15200 16643 15204
rect 16659 15260 16723 15264
rect 16659 15204 16663 15260
rect 16663 15204 16719 15260
rect 16719 15204 16723 15260
rect 16659 15200 16723 15204
rect 16739 15260 16803 15264
rect 16739 15204 16743 15260
rect 16743 15204 16799 15260
rect 16799 15204 16803 15260
rect 16739 15200 16803 15204
rect 2895 14716 2959 14720
rect 2895 14660 2899 14716
rect 2899 14660 2955 14716
rect 2955 14660 2959 14716
rect 2895 14656 2959 14660
rect 2975 14716 3039 14720
rect 2975 14660 2979 14716
rect 2979 14660 3035 14716
rect 3035 14660 3039 14716
rect 2975 14656 3039 14660
rect 3055 14716 3119 14720
rect 3055 14660 3059 14716
rect 3059 14660 3115 14716
rect 3115 14660 3119 14716
rect 3055 14656 3119 14660
rect 3135 14716 3199 14720
rect 3135 14660 3139 14716
rect 3139 14660 3195 14716
rect 3195 14660 3199 14716
rect 3135 14656 3199 14660
rect 6782 14716 6846 14720
rect 6782 14660 6786 14716
rect 6786 14660 6842 14716
rect 6842 14660 6846 14716
rect 6782 14656 6846 14660
rect 6862 14716 6926 14720
rect 6862 14660 6866 14716
rect 6866 14660 6922 14716
rect 6922 14660 6926 14716
rect 6862 14656 6926 14660
rect 6942 14716 7006 14720
rect 6942 14660 6946 14716
rect 6946 14660 7002 14716
rect 7002 14660 7006 14716
rect 6942 14656 7006 14660
rect 7022 14716 7086 14720
rect 7022 14660 7026 14716
rect 7026 14660 7082 14716
rect 7082 14660 7086 14716
rect 7022 14656 7086 14660
rect 10669 14716 10733 14720
rect 10669 14660 10673 14716
rect 10673 14660 10729 14716
rect 10729 14660 10733 14716
rect 10669 14656 10733 14660
rect 10749 14716 10813 14720
rect 10749 14660 10753 14716
rect 10753 14660 10809 14716
rect 10809 14660 10813 14716
rect 10749 14656 10813 14660
rect 10829 14716 10893 14720
rect 10829 14660 10833 14716
rect 10833 14660 10889 14716
rect 10889 14660 10893 14716
rect 10829 14656 10893 14660
rect 10909 14716 10973 14720
rect 10909 14660 10913 14716
rect 10913 14660 10969 14716
rect 10969 14660 10973 14716
rect 10909 14656 10973 14660
rect 14556 14716 14620 14720
rect 14556 14660 14560 14716
rect 14560 14660 14616 14716
rect 14616 14660 14620 14716
rect 14556 14656 14620 14660
rect 14636 14716 14700 14720
rect 14636 14660 14640 14716
rect 14640 14660 14696 14716
rect 14696 14660 14700 14716
rect 14636 14656 14700 14660
rect 14716 14716 14780 14720
rect 14716 14660 14720 14716
rect 14720 14660 14776 14716
rect 14776 14660 14780 14716
rect 14716 14656 14780 14660
rect 14796 14716 14860 14720
rect 14796 14660 14800 14716
rect 14800 14660 14856 14716
rect 14856 14660 14860 14716
rect 14796 14656 14860 14660
rect 4838 14172 4902 14176
rect 4838 14116 4842 14172
rect 4842 14116 4898 14172
rect 4898 14116 4902 14172
rect 4838 14112 4902 14116
rect 4918 14172 4982 14176
rect 4918 14116 4922 14172
rect 4922 14116 4978 14172
rect 4978 14116 4982 14172
rect 4918 14112 4982 14116
rect 4998 14172 5062 14176
rect 4998 14116 5002 14172
rect 5002 14116 5058 14172
rect 5058 14116 5062 14172
rect 4998 14112 5062 14116
rect 5078 14172 5142 14176
rect 5078 14116 5082 14172
rect 5082 14116 5138 14172
rect 5138 14116 5142 14172
rect 5078 14112 5142 14116
rect 8725 14172 8789 14176
rect 8725 14116 8729 14172
rect 8729 14116 8785 14172
rect 8785 14116 8789 14172
rect 8725 14112 8789 14116
rect 8805 14172 8869 14176
rect 8805 14116 8809 14172
rect 8809 14116 8865 14172
rect 8865 14116 8869 14172
rect 8805 14112 8869 14116
rect 8885 14172 8949 14176
rect 8885 14116 8889 14172
rect 8889 14116 8945 14172
rect 8945 14116 8949 14172
rect 8885 14112 8949 14116
rect 8965 14172 9029 14176
rect 8965 14116 8969 14172
rect 8969 14116 9025 14172
rect 9025 14116 9029 14172
rect 8965 14112 9029 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 16499 14172 16563 14176
rect 16499 14116 16503 14172
rect 16503 14116 16559 14172
rect 16559 14116 16563 14172
rect 16499 14112 16563 14116
rect 16579 14172 16643 14176
rect 16579 14116 16583 14172
rect 16583 14116 16639 14172
rect 16639 14116 16643 14172
rect 16579 14112 16643 14116
rect 16659 14172 16723 14176
rect 16659 14116 16663 14172
rect 16663 14116 16719 14172
rect 16719 14116 16723 14172
rect 16659 14112 16723 14116
rect 16739 14172 16803 14176
rect 16739 14116 16743 14172
rect 16743 14116 16799 14172
rect 16799 14116 16803 14172
rect 16739 14112 16803 14116
rect 2895 13628 2959 13632
rect 2895 13572 2899 13628
rect 2899 13572 2955 13628
rect 2955 13572 2959 13628
rect 2895 13568 2959 13572
rect 2975 13628 3039 13632
rect 2975 13572 2979 13628
rect 2979 13572 3035 13628
rect 3035 13572 3039 13628
rect 2975 13568 3039 13572
rect 3055 13628 3119 13632
rect 3055 13572 3059 13628
rect 3059 13572 3115 13628
rect 3115 13572 3119 13628
rect 3055 13568 3119 13572
rect 3135 13628 3199 13632
rect 3135 13572 3139 13628
rect 3139 13572 3195 13628
rect 3195 13572 3199 13628
rect 3135 13568 3199 13572
rect 6782 13628 6846 13632
rect 6782 13572 6786 13628
rect 6786 13572 6842 13628
rect 6842 13572 6846 13628
rect 6782 13568 6846 13572
rect 6862 13628 6926 13632
rect 6862 13572 6866 13628
rect 6866 13572 6922 13628
rect 6922 13572 6926 13628
rect 6862 13568 6926 13572
rect 6942 13628 7006 13632
rect 6942 13572 6946 13628
rect 6946 13572 7002 13628
rect 7002 13572 7006 13628
rect 6942 13568 7006 13572
rect 7022 13628 7086 13632
rect 7022 13572 7026 13628
rect 7026 13572 7082 13628
rect 7082 13572 7086 13628
rect 7022 13568 7086 13572
rect 10669 13628 10733 13632
rect 10669 13572 10673 13628
rect 10673 13572 10729 13628
rect 10729 13572 10733 13628
rect 10669 13568 10733 13572
rect 10749 13628 10813 13632
rect 10749 13572 10753 13628
rect 10753 13572 10809 13628
rect 10809 13572 10813 13628
rect 10749 13568 10813 13572
rect 10829 13628 10893 13632
rect 10829 13572 10833 13628
rect 10833 13572 10889 13628
rect 10889 13572 10893 13628
rect 10829 13568 10893 13572
rect 10909 13628 10973 13632
rect 10909 13572 10913 13628
rect 10913 13572 10969 13628
rect 10969 13572 10973 13628
rect 10909 13568 10973 13572
rect 14556 13628 14620 13632
rect 14556 13572 14560 13628
rect 14560 13572 14616 13628
rect 14616 13572 14620 13628
rect 14556 13568 14620 13572
rect 14636 13628 14700 13632
rect 14636 13572 14640 13628
rect 14640 13572 14696 13628
rect 14696 13572 14700 13628
rect 14636 13568 14700 13572
rect 14716 13628 14780 13632
rect 14716 13572 14720 13628
rect 14720 13572 14776 13628
rect 14776 13572 14780 13628
rect 14716 13568 14780 13572
rect 14796 13628 14860 13632
rect 14796 13572 14800 13628
rect 14800 13572 14856 13628
rect 14856 13572 14860 13628
rect 14796 13568 14860 13572
rect 4838 13084 4902 13088
rect 4838 13028 4842 13084
rect 4842 13028 4898 13084
rect 4898 13028 4902 13084
rect 4838 13024 4902 13028
rect 4918 13084 4982 13088
rect 4918 13028 4922 13084
rect 4922 13028 4978 13084
rect 4978 13028 4982 13084
rect 4918 13024 4982 13028
rect 4998 13084 5062 13088
rect 4998 13028 5002 13084
rect 5002 13028 5058 13084
rect 5058 13028 5062 13084
rect 4998 13024 5062 13028
rect 5078 13084 5142 13088
rect 5078 13028 5082 13084
rect 5082 13028 5138 13084
rect 5138 13028 5142 13084
rect 5078 13024 5142 13028
rect 8725 13084 8789 13088
rect 8725 13028 8729 13084
rect 8729 13028 8785 13084
rect 8785 13028 8789 13084
rect 8725 13024 8789 13028
rect 8805 13084 8869 13088
rect 8805 13028 8809 13084
rect 8809 13028 8865 13084
rect 8865 13028 8869 13084
rect 8805 13024 8869 13028
rect 8885 13084 8949 13088
rect 8885 13028 8889 13084
rect 8889 13028 8945 13084
rect 8945 13028 8949 13084
rect 8885 13024 8949 13028
rect 8965 13084 9029 13088
rect 8965 13028 8969 13084
rect 8969 13028 9025 13084
rect 9025 13028 9029 13084
rect 8965 13024 9029 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 16499 13084 16563 13088
rect 16499 13028 16503 13084
rect 16503 13028 16559 13084
rect 16559 13028 16563 13084
rect 16499 13024 16563 13028
rect 16579 13084 16643 13088
rect 16579 13028 16583 13084
rect 16583 13028 16639 13084
rect 16639 13028 16643 13084
rect 16579 13024 16643 13028
rect 16659 13084 16723 13088
rect 16659 13028 16663 13084
rect 16663 13028 16719 13084
rect 16719 13028 16723 13084
rect 16659 13024 16723 13028
rect 16739 13084 16803 13088
rect 16739 13028 16743 13084
rect 16743 13028 16799 13084
rect 16799 13028 16803 13084
rect 16739 13024 16803 13028
rect 2895 12540 2959 12544
rect 2895 12484 2899 12540
rect 2899 12484 2955 12540
rect 2955 12484 2959 12540
rect 2895 12480 2959 12484
rect 2975 12540 3039 12544
rect 2975 12484 2979 12540
rect 2979 12484 3035 12540
rect 3035 12484 3039 12540
rect 2975 12480 3039 12484
rect 3055 12540 3119 12544
rect 3055 12484 3059 12540
rect 3059 12484 3115 12540
rect 3115 12484 3119 12540
rect 3055 12480 3119 12484
rect 3135 12540 3199 12544
rect 3135 12484 3139 12540
rect 3139 12484 3195 12540
rect 3195 12484 3199 12540
rect 3135 12480 3199 12484
rect 6782 12540 6846 12544
rect 6782 12484 6786 12540
rect 6786 12484 6842 12540
rect 6842 12484 6846 12540
rect 6782 12480 6846 12484
rect 6862 12540 6926 12544
rect 6862 12484 6866 12540
rect 6866 12484 6922 12540
rect 6922 12484 6926 12540
rect 6862 12480 6926 12484
rect 6942 12540 7006 12544
rect 6942 12484 6946 12540
rect 6946 12484 7002 12540
rect 7002 12484 7006 12540
rect 6942 12480 7006 12484
rect 7022 12540 7086 12544
rect 7022 12484 7026 12540
rect 7026 12484 7082 12540
rect 7082 12484 7086 12540
rect 7022 12480 7086 12484
rect 10669 12540 10733 12544
rect 10669 12484 10673 12540
rect 10673 12484 10729 12540
rect 10729 12484 10733 12540
rect 10669 12480 10733 12484
rect 10749 12540 10813 12544
rect 10749 12484 10753 12540
rect 10753 12484 10809 12540
rect 10809 12484 10813 12540
rect 10749 12480 10813 12484
rect 10829 12540 10893 12544
rect 10829 12484 10833 12540
rect 10833 12484 10889 12540
rect 10889 12484 10893 12540
rect 10829 12480 10893 12484
rect 10909 12540 10973 12544
rect 10909 12484 10913 12540
rect 10913 12484 10969 12540
rect 10969 12484 10973 12540
rect 10909 12480 10973 12484
rect 14556 12540 14620 12544
rect 14556 12484 14560 12540
rect 14560 12484 14616 12540
rect 14616 12484 14620 12540
rect 14556 12480 14620 12484
rect 14636 12540 14700 12544
rect 14636 12484 14640 12540
rect 14640 12484 14696 12540
rect 14696 12484 14700 12540
rect 14636 12480 14700 12484
rect 14716 12540 14780 12544
rect 14716 12484 14720 12540
rect 14720 12484 14776 12540
rect 14776 12484 14780 12540
rect 14716 12480 14780 12484
rect 14796 12540 14860 12544
rect 14796 12484 14800 12540
rect 14800 12484 14856 12540
rect 14856 12484 14860 12540
rect 14796 12480 14860 12484
rect 4838 11996 4902 12000
rect 4838 11940 4842 11996
rect 4842 11940 4898 11996
rect 4898 11940 4902 11996
rect 4838 11936 4902 11940
rect 4918 11996 4982 12000
rect 4918 11940 4922 11996
rect 4922 11940 4978 11996
rect 4978 11940 4982 11996
rect 4918 11936 4982 11940
rect 4998 11996 5062 12000
rect 4998 11940 5002 11996
rect 5002 11940 5058 11996
rect 5058 11940 5062 11996
rect 4998 11936 5062 11940
rect 5078 11996 5142 12000
rect 5078 11940 5082 11996
rect 5082 11940 5138 11996
rect 5138 11940 5142 11996
rect 5078 11936 5142 11940
rect 8725 11996 8789 12000
rect 8725 11940 8729 11996
rect 8729 11940 8785 11996
rect 8785 11940 8789 11996
rect 8725 11936 8789 11940
rect 8805 11996 8869 12000
rect 8805 11940 8809 11996
rect 8809 11940 8865 11996
rect 8865 11940 8869 11996
rect 8805 11936 8869 11940
rect 8885 11996 8949 12000
rect 8885 11940 8889 11996
rect 8889 11940 8945 11996
rect 8945 11940 8949 11996
rect 8885 11936 8949 11940
rect 8965 11996 9029 12000
rect 8965 11940 8969 11996
rect 8969 11940 9025 11996
rect 9025 11940 9029 11996
rect 8965 11936 9029 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 16499 11996 16563 12000
rect 16499 11940 16503 11996
rect 16503 11940 16559 11996
rect 16559 11940 16563 11996
rect 16499 11936 16563 11940
rect 16579 11996 16643 12000
rect 16579 11940 16583 11996
rect 16583 11940 16639 11996
rect 16639 11940 16643 11996
rect 16579 11936 16643 11940
rect 16659 11996 16723 12000
rect 16659 11940 16663 11996
rect 16663 11940 16719 11996
rect 16719 11940 16723 11996
rect 16659 11936 16723 11940
rect 16739 11996 16803 12000
rect 16739 11940 16743 11996
rect 16743 11940 16799 11996
rect 16799 11940 16803 11996
rect 16739 11936 16803 11940
rect 2895 11452 2959 11456
rect 2895 11396 2899 11452
rect 2899 11396 2955 11452
rect 2955 11396 2959 11452
rect 2895 11392 2959 11396
rect 2975 11452 3039 11456
rect 2975 11396 2979 11452
rect 2979 11396 3035 11452
rect 3035 11396 3039 11452
rect 2975 11392 3039 11396
rect 3055 11452 3119 11456
rect 3055 11396 3059 11452
rect 3059 11396 3115 11452
rect 3115 11396 3119 11452
rect 3055 11392 3119 11396
rect 3135 11452 3199 11456
rect 3135 11396 3139 11452
rect 3139 11396 3195 11452
rect 3195 11396 3199 11452
rect 3135 11392 3199 11396
rect 6782 11452 6846 11456
rect 6782 11396 6786 11452
rect 6786 11396 6842 11452
rect 6842 11396 6846 11452
rect 6782 11392 6846 11396
rect 6862 11452 6926 11456
rect 6862 11396 6866 11452
rect 6866 11396 6922 11452
rect 6922 11396 6926 11452
rect 6862 11392 6926 11396
rect 6942 11452 7006 11456
rect 6942 11396 6946 11452
rect 6946 11396 7002 11452
rect 7002 11396 7006 11452
rect 6942 11392 7006 11396
rect 7022 11452 7086 11456
rect 7022 11396 7026 11452
rect 7026 11396 7082 11452
rect 7082 11396 7086 11452
rect 7022 11392 7086 11396
rect 10669 11452 10733 11456
rect 10669 11396 10673 11452
rect 10673 11396 10729 11452
rect 10729 11396 10733 11452
rect 10669 11392 10733 11396
rect 10749 11452 10813 11456
rect 10749 11396 10753 11452
rect 10753 11396 10809 11452
rect 10809 11396 10813 11452
rect 10749 11392 10813 11396
rect 10829 11452 10893 11456
rect 10829 11396 10833 11452
rect 10833 11396 10889 11452
rect 10889 11396 10893 11452
rect 10829 11392 10893 11396
rect 10909 11452 10973 11456
rect 10909 11396 10913 11452
rect 10913 11396 10969 11452
rect 10969 11396 10973 11452
rect 10909 11392 10973 11396
rect 14556 11452 14620 11456
rect 14556 11396 14560 11452
rect 14560 11396 14616 11452
rect 14616 11396 14620 11452
rect 14556 11392 14620 11396
rect 14636 11452 14700 11456
rect 14636 11396 14640 11452
rect 14640 11396 14696 11452
rect 14696 11396 14700 11452
rect 14636 11392 14700 11396
rect 14716 11452 14780 11456
rect 14716 11396 14720 11452
rect 14720 11396 14776 11452
rect 14776 11396 14780 11452
rect 14716 11392 14780 11396
rect 14796 11452 14860 11456
rect 14796 11396 14800 11452
rect 14800 11396 14856 11452
rect 14856 11396 14860 11452
rect 14796 11392 14860 11396
rect 4838 10908 4902 10912
rect 4838 10852 4842 10908
rect 4842 10852 4898 10908
rect 4898 10852 4902 10908
rect 4838 10848 4902 10852
rect 4918 10908 4982 10912
rect 4918 10852 4922 10908
rect 4922 10852 4978 10908
rect 4978 10852 4982 10908
rect 4918 10848 4982 10852
rect 4998 10908 5062 10912
rect 4998 10852 5002 10908
rect 5002 10852 5058 10908
rect 5058 10852 5062 10908
rect 4998 10848 5062 10852
rect 5078 10908 5142 10912
rect 5078 10852 5082 10908
rect 5082 10852 5138 10908
rect 5138 10852 5142 10908
rect 5078 10848 5142 10852
rect 8725 10908 8789 10912
rect 8725 10852 8729 10908
rect 8729 10852 8785 10908
rect 8785 10852 8789 10908
rect 8725 10848 8789 10852
rect 8805 10908 8869 10912
rect 8805 10852 8809 10908
rect 8809 10852 8865 10908
rect 8865 10852 8869 10908
rect 8805 10848 8869 10852
rect 8885 10908 8949 10912
rect 8885 10852 8889 10908
rect 8889 10852 8945 10908
rect 8945 10852 8949 10908
rect 8885 10848 8949 10852
rect 8965 10908 9029 10912
rect 8965 10852 8969 10908
rect 8969 10852 9025 10908
rect 9025 10852 9029 10908
rect 8965 10848 9029 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 16499 10908 16563 10912
rect 16499 10852 16503 10908
rect 16503 10852 16559 10908
rect 16559 10852 16563 10908
rect 16499 10848 16563 10852
rect 16579 10908 16643 10912
rect 16579 10852 16583 10908
rect 16583 10852 16639 10908
rect 16639 10852 16643 10908
rect 16579 10848 16643 10852
rect 16659 10908 16723 10912
rect 16659 10852 16663 10908
rect 16663 10852 16719 10908
rect 16719 10852 16723 10908
rect 16659 10848 16723 10852
rect 16739 10908 16803 10912
rect 16739 10852 16743 10908
rect 16743 10852 16799 10908
rect 16799 10852 16803 10908
rect 16739 10848 16803 10852
rect 2895 10364 2959 10368
rect 2895 10308 2899 10364
rect 2899 10308 2955 10364
rect 2955 10308 2959 10364
rect 2895 10304 2959 10308
rect 2975 10364 3039 10368
rect 2975 10308 2979 10364
rect 2979 10308 3035 10364
rect 3035 10308 3039 10364
rect 2975 10304 3039 10308
rect 3055 10364 3119 10368
rect 3055 10308 3059 10364
rect 3059 10308 3115 10364
rect 3115 10308 3119 10364
rect 3055 10304 3119 10308
rect 3135 10364 3199 10368
rect 3135 10308 3139 10364
rect 3139 10308 3195 10364
rect 3195 10308 3199 10364
rect 3135 10304 3199 10308
rect 6782 10364 6846 10368
rect 6782 10308 6786 10364
rect 6786 10308 6842 10364
rect 6842 10308 6846 10364
rect 6782 10304 6846 10308
rect 6862 10364 6926 10368
rect 6862 10308 6866 10364
rect 6866 10308 6922 10364
rect 6922 10308 6926 10364
rect 6862 10304 6926 10308
rect 6942 10364 7006 10368
rect 6942 10308 6946 10364
rect 6946 10308 7002 10364
rect 7002 10308 7006 10364
rect 6942 10304 7006 10308
rect 7022 10364 7086 10368
rect 7022 10308 7026 10364
rect 7026 10308 7082 10364
rect 7082 10308 7086 10364
rect 7022 10304 7086 10308
rect 10669 10364 10733 10368
rect 10669 10308 10673 10364
rect 10673 10308 10729 10364
rect 10729 10308 10733 10364
rect 10669 10304 10733 10308
rect 10749 10364 10813 10368
rect 10749 10308 10753 10364
rect 10753 10308 10809 10364
rect 10809 10308 10813 10364
rect 10749 10304 10813 10308
rect 10829 10364 10893 10368
rect 10829 10308 10833 10364
rect 10833 10308 10889 10364
rect 10889 10308 10893 10364
rect 10829 10304 10893 10308
rect 10909 10364 10973 10368
rect 10909 10308 10913 10364
rect 10913 10308 10969 10364
rect 10969 10308 10973 10364
rect 10909 10304 10973 10308
rect 14556 10364 14620 10368
rect 14556 10308 14560 10364
rect 14560 10308 14616 10364
rect 14616 10308 14620 10364
rect 14556 10304 14620 10308
rect 14636 10364 14700 10368
rect 14636 10308 14640 10364
rect 14640 10308 14696 10364
rect 14696 10308 14700 10364
rect 14636 10304 14700 10308
rect 14716 10364 14780 10368
rect 14716 10308 14720 10364
rect 14720 10308 14776 10364
rect 14776 10308 14780 10364
rect 14716 10304 14780 10308
rect 14796 10364 14860 10368
rect 14796 10308 14800 10364
rect 14800 10308 14856 10364
rect 14856 10308 14860 10364
rect 14796 10304 14860 10308
rect 4838 9820 4902 9824
rect 4838 9764 4842 9820
rect 4842 9764 4898 9820
rect 4898 9764 4902 9820
rect 4838 9760 4902 9764
rect 4918 9820 4982 9824
rect 4918 9764 4922 9820
rect 4922 9764 4978 9820
rect 4978 9764 4982 9820
rect 4918 9760 4982 9764
rect 4998 9820 5062 9824
rect 4998 9764 5002 9820
rect 5002 9764 5058 9820
rect 5058 9764 5062 9820
rect 4998 9760 5062 9764
rect 5078 9820 5142 9824
rect 5078 9764 5082 9820
rect 5082 9764 5138 9820
rect 5138 9764 5142 9820
rect 5078 9760 5142 9764
rect 8725 9820 8789 9824
rect 8725 9764 8729 9820
rect 8729 9764 8785 9820
rect 8785 9764 8789 9820
rect 8725 9760 8789 9764
rect 8805 9820 8869 9824
rect 8805 9764 8809 9820
rect 8809 9764 8865 9820
rect 8865 9764 8869 9820
rect 8805 9760 8869 9764
rect 8885 9820 8949 9824
rect 8885 9764 8889 9820
rect 8889 9764 8945 9820
rect 8945 9764 8949 9820
rect 8885 9760 8949 9764
rect 8965 9820 9029 9824
rect 8965 9764 8969 9820
rect 8969 9764 9025 9820
rect 9025 9764 9029 9820
rect 8965 9760 9029 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 16499 9820 16563 9824
rect 16499 9764 16503 9820
rect 16503 9764 16559 9820
rect 16559 9764 16563 9820
rect 16499 9760 16563 9764
rect 16579 9820 16643 9824
rect 16579 9764 16583 9820
rect 16583 9764 16639 9820
rect 16639 9764 16643 9820
rect 16579 9760 16643 9764
rect 16659 9820 16723 9824
rect 16659 9764 16663 9820
rect 16663 9764 16719 9820
rect 16719 9764 16723 9820
rect 16659 9760 16723 9764
rect 16739 9820 16803 9824
rect 16739 9764 16743 9820
rect 16743 9764 16799 9820
rect 16799 9764 16803 9820
rect 16739 9760 16803 9764
rect 2895 9276 2959 9280
rect 2895 9220 2899 9276
rect 2899 9220 2955 9276
rect 2955 9220 2959 9276
rect 2895 9216 2959 9220
rect 2975 9276 3039 9280
rect 2975 9220 2979 9276
rect 2979 9220 3035 9276
rect 3035 9220 3039 9276
rect 2975 9216 3039 9220
rect 3055 9276 3119 9280
rect 3055 9220 3059 9276
rect 3059 9220 3115 9276
rect 3115 9220 3119 9276
rect 3055 9216 3119 9220
rect 3135 9276 3199 9280
rect 3135 9220 3139 9276
rect 3139 9220 3195 9276
rect 3195 9220 3199 9276
rect 3135 9216 3199 9220
rect 6782 9276 6846 9280
rect 6782 9220 6786 9276
rect 6786 9220 6842 9276
rect 6842 9220 6846 9276
rect 6782 9216 6846 9220
rect 6862 9276 6926 9280
rect 6862 9220 6866 9276
rect 6866 9220 6922 9276
rect 6922 9220 6926 9276
rect 6862 9216 6926 9220
rect 6942 9276 7006 9280
rect 6942 9220 6946 9276
rect 6946 9220 7002 9276
rect 7002 9220 7006 9276
rect 6942 9216 7006 9220
rect 7022 9276 7086 9280
rect 7022 9220 7026 9276
rect 7026 9220 7082 9276
rect 7082 9220 7086 9276
rect 7022 9216 7086 9220
rect 10669 9276 10733 9280
rect 10669 9220 10673 9276
rect 10673 9220 10729 9276
rect 10729 9220 10733 9276
rect 10669 9216 10733 9220
rect 10749 9276 10813 9280
rect 10749 9220 10753 9276
rect 10753 9220 10809 9276
rect 10809 9220 10813 9276
rect 10749 9216 10813 9220
rect 10829 9276 10893 9280
rect 10829 9220 10833 9276
rect 10833 9220 10889 9276
rect 10889 9220 10893 9276
rect 10829 9216 10893 9220
rect 10909 9276 10973 9280
rect 10909 9220 10913 9276
rect 10913 9220 10969 9276
rect 10969 9220 10973 9276
rect 10909 9216 10973 9220
rect 14556 9276 14620 9280
rect 14556 9220 14560 9276
rect 14560 9220 14616 9276
rect 14616 9220 14620 9276
rect 14556 9216 14620 9220
rect 14636 9276 14700 9280
rect 14636 9220 14640 9276
rect 14640 9220 14696 9276
rect 14696 9220 14700 9276
rect 14636 9216 14700 9220
rect 14716 9276 14780 9280
rect 14716 9220 14720 9276
rect 14720 9220 14776 9276
rect 14776 9220 14780 9276
rect 14716 9216 14780 9220
rect 14796 9276 14860 9280
rect 14796 9220 14800 9276
rect 14800 9220 14856 9276
rect 14856 9220 14860 9276
rect 14796 9216 14860 9220
rect 4838 8732 4902 8736
rect 4838 8676 4842 8732
rect 4842 8676 4898 8732
rect 4898 8676 4902 8732
rect 4838 8672 4902 8676
rect 4918 8732 4982 8736
rect 4918 8676 4922 8732
rect 4922 8676 4978 8732
rect 4978 8676 4982 8732
rect 4918 8672 4982 8676
rect 4998 8732 5062 8736
rect 4998 8676 5002 8732
rect 5002 8676 5058 8732
rect 5058 8676 5062 8732
rect 4998 8672 5062 8676
rect 5078 8732 5142 8736
rect 5078 8676 5082 8732
rect 5082 8676 5138 8732
rect 5138 8676 5142 8732
rect 5078 8672 5142 8676
rect 8725 8732 8789 8736
rect 8725 8676 8729 8732
rect 8729 8676 8785 8732
rect 8785 8676 8789 8732
rect 8725 8672 8789 8676
rect 8805 8732 8869 8736
rect 8805 8676 8809 8732
rect 8809 8676 8865 8732
rect 8865 8676 8869 8732
rect 8805 8672 8869 8676
rect 8885 8732 8949 8736
rect 8885 8676 8889 8732
rect 8889 8676 8945 8732
rect 8945 8676 8949 8732
rect 8885 8672 8949 8676
rect 8965 8732 9029 8736
rect 8965 8676 8969 8732
rect 8969 8676 9025 8732
rect 9025 8676 9029 8732
rect 8965 8672 9029 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 16499 8732 16563 8736
rect 16499 8676 16503 8732
rect 16503 8676 16559 8732
rect 16559 8676 16563 8732
rect 16499 8672 16563 8676
rect 16579 8732 16643 8736
rect 16579 8676 16583 8732
rect 16583 8676 16639 8732
rect 16639 8676 16643 8732
rect 16579 8672 16643 8676
rect 16659 8732 16723 8736
rect 16659 8676 16663 8732
rect 16663 8676 16719 8732
rect 16719 8676 16723 8732
rect 16659 8672 16723 8676
rect 16739 8732 16803 8736
rect 16739 8676 16743 8732
rect 16743 8676 16799 8732
rect 16799 8676 16803 8732
rect 16739 8672 16803 8676
rect 2895 8188 2959 8192
rect 2895 8132 2899 8188
rect 2899 8132 2955 8188
rect 2955 8132 2959 8188
rect 2895 8128 2959 8132
rect 2975 8188 3039 8192
rect 2975 8132 2979 8188
rect 2979 8132 3035 8188
rect 3035 8132 3039 8188
rect 2975 8128 3039 8132
rect 3055 8188 3119 8192
rect 3055 8132 3059 8188
rect 3059 8132 3115 8188
rect 3115 8132 3119 8188
rect 3055 8128 3119 8132
rect 3135 8188 3199 8192
rect 3135 8132 3139 8188
rect 3139 8132 3195 8188
rect 3195 8132 3199 8188
rect 3135 8128 3199 8132
rect 6782 8188 6846 8192
rect 6782 8132 6786 8188
rect 6786 8132 6842 8188
rect 6842 8132 6846 8188
rect 6782 8128 6846 8132
rect 6862 8188 6926 8192
rect 6862 8132 6866 8188
rect 6866 8132 6922 8188
rect 6922 8132 6926 8188
rect 6862 8128 6926 8132
rect 6942 8188 7006 8192
rect 6942 8132 6946 8188
rect 6946 8132 7002 8188
rect 7002 8132 7006 8188
rect 6942 8128 7006 8132
rect 7022 8188 7086 8192
rect 7022 8132 7026 8188
rect 7026 8132 7082 8188
rect 7082 8132 7086 8188
rect 7022 8128 7086 8132
rect 10669 8188 10733 8192
rect 10669 8132 10673 8188
rect 10673 8132 10729 8188
rect 10729 8132 10733 8188
rect 10669 8128 10733 8132
rect 10749 8188 10813 8192
rect 10749 8132 10753 8188
rect 10753 8132 10809 8188
rect 10809 8132 10813 8188
rect 10749 8128 10813 8132
rect 10829 8188 10893 8192
rect 10829 8132 10833 8188
rect 10833 8132 10889 8188
rect 10889 8132 10893 8188
rect 10829 8128 10893 8132
rect 10909 8188 10973 8192
rect 10909 8132 10913 8188
rect 10913 8132 10969 8188
rect 10969 8132 10973 8188
rect 10909 8128 10973 8132
rect 14556 8188 14620 8192
rect 14556 8132 14560 8188
rect 14560 8132 14616 8188
rect 14616 8132 14620 8188
rect 14556 8128 14620 8132
rect 14636 8188 14700 8192
rect 14636 8132 14640 8188
rect 14640 8132 14696 8188
rect 14696 8132 14700 8188
rect 14636 8128 14700 8132
rect 14716 8188 14780 8192
rect 14716 8132 14720 8188
rect 14720 8132 14776 8188
rect 14776 8132 14780 8188
rect 14716 8128 14780 8132
rect 14796 8188 14860 8192
rect 14796 8132 14800 8188
rect 14800 8132 14856 8188
rect 14856 8132 14860 8188
rect 14796 8128 14860 8132
rect 4838 7644 4902 7648
rect 4838 7588 4842 7644
rect 4842 7588 4898 7644
rect 4898 7588 4902 7644
rect 4838 7584 4902 7588
rect 4918 7644 4982 7648
rect 4918 7588 4922 7644
rect 4922 7588 4978 7644
rect 4978 7588 4982 7644
rect 4918 7584 4982 7588
rect 4998 7644 5062 7648
rect 4998 7588 5002 7644
rect 5002 7588 5058 7644
rect 5058 7588 5062 7644
rect 4998 7584 5062 7588
rect 5078 7644 5142 7648
rect 5078 7588 5082 7644
rect 5082 7588 5138 7644
rect 5138 7588 5142 7644
rect 5078 7584 5142 7588
rect 8725 7644 8789 7648
rect 8725 7588 8729 7644
rect 8729 7588 8785 7644
rect 8785 7588 8789 7644
rect 8725 7584 8789 7588
rect 8805 7644 8869 7648
rect 8805 7588 8809 7644
rect 8809 7588 8865 7644
rect 8865 7588 8869 7644
rect 8805 7584 8869 7588
rect 8885 7644 8949 7648
rect 8885 7588 8889 7644
rect 8889 7588 8945 7644
rect 8945 7588 8949 7644
rect 8885 7584 8949 7588
rect 8965 7644 9029 7648
rect 8965 7588 8969 7644
rect 8969 7588 9025 7644
rect 9025 7588 9029 7644
rect 8965 7584 9029 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 16499 7644 16563 7648
rect 16499 7588 16503 7644
rect 16503 7588 16559 7644
rect 16559 7588 16563 7644
rect 16499 7584 16563 7588
rect 16579 7644 16643 7648
rect 16579 7588 16583 7644
rect 16583 7588 16639 7644
rect 16639 7588 16643 7644
rect 16579 7584 16643 7588
rect 16659 7644 16723 7648
rect 16659 7588 16663 7644
rect 16663 7588 16719 7644
rect 16719 7588 16723 7644
rect 16659 7584 16723 7588
rect 16739 7644 16803 7648
rect 16739 7588 16743 7644
rect 16743 7588 16799 7644
rect 16799 7588 16803 7644
rect 16739 7584 16803 7588
rect 2895 7100 2959 7104
rect 2895 7044 2899 7100
rect 2899 7044 2955 7100
rect 2955 7044 2959 7100
rect 2895 7040 2959 7044
rect 2975 7100 3039 7104
rect 2975 7044 2979 7100
rect 2979 7044 3035 7100
rect 3035 7044 3039 7100
rect 2975 7040 3039 7044
rect 3055 7100 3119 7104
rect 3055 7044 3059 7100
rect 3059 7044 3115 7100
rect 3115 7044 3119 7100
rect 3055 7040 3119 7044
rect 3135 7100 3199 7104
rect 3135 7044 3139 7100
rect 3139 7044 3195 7100
rect 3195 7044 3199 7100
rect 3135 7040 3199 7044
rect 6782 7100 6846 7104
rect 6782 7044 6786 7100
rect 6786 7044 6842 7100
rect 6842 7044 6846 7100
rect 6782 7040 6846 7044
rect 6862 7100 6926 7104
rect 6862 7044 6866 7100
rect 6866 7044 6922 7100
rect 6922 7044 6926 7100
rect 6862 7040 6926 7044
rect 6942 7100 7006 7104
rect 6942 7044 6946 7100
rect 6946 7044 7002 7100
rect 7002 7044 7006 7100
rect 6942 7040 7006 7044
rect 7022 7100 7086 7104
rect 7022 7044 7026 7100
rect 7026 7044 7082 7100
rect 7082 7044 7086 7100
rect 7022 7040 7086 7044
rect 10669 7100 10733 7104
rect 10669 7044 10673 7100
rect 10673 7044 10729 7100
rect 10729 7044 10733 7100
rect 10669 7040 10733 7044
rect 10749 7100 10813 7104
rect 10749 7044 10753 7100
rect 10753 7044 10809 7100
rect 10809 7044 10813 7100
rect 10749 7040 10813 7044
rect 10829 7100 10893 7104
rect 10829 7044 10833 7100
rect 10833 7044 10889 7100
rect 10889 7044 10893 7100
rect 10829 7040 10893 7044
rect 10909 7100 10973 7104
rect 10909 7044 10913 7100
rect 10913 7044 10969 7100
rect 10969 7044 10973 7100
rect 10909 7040 10973 7044
rect 14556 7100 14620 7104
rect 14556 7044 14560 7100
rect 14560 7044 14616 7100
rect 14616 7044 14620 7100
rect 14556 7040 14620 7044
rect 14636 7100 14700 7104
rect 14636 7044 14640 7100
rect 14640 7044 14696 7100
rect 14696 7044 14700 7100
rect 14636 7040 14700 7044
rect 14716 7100 14780 7104
rect 14716 7044 14720 7100
rect 14720 7044 14776 7100
rect 14776 7044 14780 7100
rect 14716 7040 14780 7044
rect 14796 7100 14860 7104
rect 14796 7044 14800 7100
rect 14800 7044 14856 7100
rect 14856 7044 14860 7100
rect 14796 7040 14860 7044
rect 4838 6556 4902 6560
rect 4838 6500 4842 6556
rect 4842 6500 4898 6556
rect 4898 6500 4902 6556
rect 4838 6496 4902 6500
rect 4918 6556 4982 6560
rect 4918 6500 4922 6556
rect 4922 6500 4978 6556
rect 4978 6500 4982 6556
rect 4918 6496 4982 6500
rect 4998 6556 5062 6560
rect 4998 6500 5002 6556
rect 5002 6500 5058 6556
rect 5058 6500 5062 6556
rect 4998 6496 5062 6500
rect 5078 6556 5142 6560
rect 5078 6500 5082 6556
rect 5082 6500 5138 6556
rect 5138 6500 5142 6556
rect 5078 6496 5142 6500
rect 8725 6556 8789 6560
rect 8725 6500 8729 6556
rect 8729 6500 8785 6556
rect 8785 6500 8789 6556
rect 8725 6496 8789 6500
rect 8805 6556 8869 6560
rect 8805 6500 8809 6556
rect 8809 6500 8865 6556
rect 8865 6500 8869 6556
rect 8805 6496 8869 6500
rect 8885 6556 8949 6560
rect 8885 6500 8889 6556
rect 8889 6500 8945 6556
rect 8945 6500 8949 6556
rect 8885 6496 8949 6500
rect 8965 6556 9029 6560
rect 8965 6500 8969 6556
rect 8969 6500 9025 6556
rect 9025 6500 9029 6556
rect 8965 6496 9029 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 16499 6556 16563 6560
rect 16499 6500 16503 6556
rect 16503 6500 16559 6556
rect 16559 6500 16563 6556
rect 16499 6496 16563 6500
rect 16579 6556 16643 6560
rect 16579 6500 16583 6556
rect 16583 6500 16639 6556
rect 16639 6500 16643 6556
rect 16579 6496 16643 6500
rect 16659 6556 16723 6560
rect 16659 6500 16663 6556
rect 16663 6500 16719 6556
rect 16719 6500 16723 6556
rect 16659 6496 16723 6500
rect 16739 6556 16803 6560
rect 16739 6500 16743 6556
rect 16743 6500 16799 6556
rect 16799 6500 16803 6556
rect 16739 6496 16803 6500
rect 2895 6012 2959 6016
rect 2895 5956 2899 6012
rect 2899 5956 2955 6012
rect 2955 5956 2959 6012
rect 2895 5952 2959 5956
rect 2975 6012 3039 6016
rect 2975 5956 2979 6012
rect 2979 5956 3035 6012
rect 3035 5956 3039 6012
rect 2975 5952 3039 5956
rect 3055 6012 3119 6016
rect 3055 5956 3059 6012
rect 3059 5956 3115 6012
rect 3115 5956 3119 6012
rect 3055 5952 3119 5956
rect 3135 6012 3199 6016
rect 3135 5956 3139 6012
rect 3139 5956 3195 6012
rect 3195 5956 3199 6012
rect 3135 5952 3199 5956
rect 6782 6012 6846 6016
rect 6782 5956 6786 6012
rect 6786 5956 6842 6012
rect 6842 5956 6846 6012
rect 6782 5952 6846 5956
rect 6862 6012 6926 6016
rect 6862 5956 6866 6012
rect 6866 5956 6922 6012
rect 6922 5956 6926 6012
rect 6862 5952 6926 5956
rect 6942 6012 7006 6016
rect 6942 5956 6946 6012
rect 6946 5956 7002 6012
rect 7002 5956 7006 6012
rect 6942 5952 7006 5956
rect 7022 6012 7086 6016
rect 7022 5956 7026 6012
rect 7026 5956 7082 6012
rect 7082 5956 7086 6012
rect 7022 5952 7086 5956
rect 10669 6012 10733 6016
rect 10669 5956 10673 6012
rect 10673 5956 10729 6012
rect 10729 5956 10733 6012
rect 10669 5952 10733 5956
rect 10749 6012 10813 6016
rect 10749 5956 10753 6012
rect 10753 5956 10809 6012
rect 10809 5956 10813 6012
rect 10749 5952 10813 5956
rect 10829 6012 10893 6016
rect 10829 5956 10833 6012
rect 10833 5956 10889 6012
rect 10889 5956 10893 6012
rect 10829 5952 10893 5956
rect 10909 6012 10973 6016
rect 10909 5956 10913 6012
rect 10913 5956 10969 6012
rect 10969 5956 10973 6012
rect 10909 5952 10973 5956
rect 14556 6012 14620 6016
rect 14556 5956 14560 6012
rect 14560 5956 14616 6012
rect 14616 5956 14620 6012
rect 14556 5952 14620 5956
rect 14636 6012 14700 6016
rect 14636 5956 14640 6012
rect 14640 5956 14696 6012
rect 14696 5956 14700 6012
rect 14636 5952 14700 5956
rect 14716 6012 14780 6016
rect 14716 5956 14720 6012
rect 14720 5956 14776 6012
rect 14776 5956 14780 6012
rect 14716 5952 14780 5956
rect 14796 6012 14860 6016
rect 14796 5956 14800 6012
rect 14800 5956 14856 6012
rect 14856 5956 14860 6012
rect 14796 5952 14860 5956
rect 4838 5468 4902 5472
rect 4838 5412 4842 5468
rect 4842 5412 4898 5468
rect 4898 5412 4902 5468
rect 4838 5408 4902 5412
rect 4918 5468 4982 5472
rect 4918 5412 4922 5468
rect 4922 5412 4978 5468
rect 4978 5412 4982 5468
rect 4918 5408 4982 5412
rect 4998 5468 5062 5472
rect 4998 5412 5002 5468
rect 5002 5412 5058 5468
rect 5058 5412 5062 5468
rect 4998 5408 5062 5412
rect 5078 5468 5142 5472
rect 5078 5412 5082 5468
rect 5082 5412 5138 5468
rect 5138 5412 5142 5468
rect 5078 5408 5142 5412
rect 8725 5468 8789 5472
rect 8725 5412 8729 5468
rect 8729 5412 8785 5468
rect 8785 5412 8789 5468
rect 8725 5408 8789 5412
rect 8805 5468 8869 5472
rect 8805 5412 8809 5468
rect 8809 5412 8865 5468
rect 8865 5412 8869 5468
rect 8805 5408 8869 5412
rect 8885 5468 8949 5472
rect 8885 5412 8889 5468
rect 8889 5412 8945 5468
rect 8945 5412 8949 5468
rect 8885 5408 8949 5412
rect 8965 5468 9029 5472
rect 8965 5412 8969 5468
rect 8969 5412 9025 5468
rect 9025 5412 9029 5468
rect 8965 5408 9029 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 16499 5468 16563 5472
rect 16499 5412 16503 5468
rect 16503 5412 16559 5468
rect 16559 5412 16563 5468
rect 16499 5408 16563 5412
rect 16579 5468 16643 5472
rect 16579 5412 16583 5468
rect 16583 5412 16639 5468
rect 16639 5412 16643 5468
rect 16579 5408 16643 5412
rect 16659 5468 16723 5472
rect 16659 5412 16663 5468
rect 16663 5412 16719 5468
rect 16719 5412 16723 5468
rect 16659 5408 16723 5412
rect 16739 5468 16803 5472
rect 16739 5412 16743 5468
rect 16743 5412 16799 5468
rect 16799 5412 16803 5468
rect 16739 5408 16803 5412
rect 2895 4924 2959 4928
rect 2895 4868 2899 4924
rect 2899 4868 2955 4924
rect 2955 4868 2959 4924
rect 2895 4864 2959 4868
rect 2975 4924 3039 4928
rect 2975 4868 2979 4924
rect 2979 4868 3035 4924
rect 3035 4868 3039 4924
rect 2975 4864 3039 4868
rect 3055 4924 3119 4928
rect 3055 4868 3059 4924
rect 3059 4868 3115 4924
rect 3115 4868 3119 4924
rect 3055 4864 3119 4868
rect 3135 4924 3199 4928
rect 3135 4868 3139 4924
rect 3139 4868 3195 4924
rect 3195 4868 3199 4924
rect 3135 4864 3199 4868
rect 6782 4924 6846 4928
rect 6782 4868 6786 4924
rect 6786 4868 6842 4924
rect 6842 4868 6846 4924
rect 6782 4864 6846 4868
rect 6862 4924 6926 4928
rect 6862 4868 6866 4924
rect 6866 4868 6922 4924
rect 6922 4868 6926 4924
rect 6862 4864 6926 4868
rect 6942 4924 7006 4928
rect 6942 4868 6946 4924
rect 6946 4868 7002 4924
rect 7002 4868 7006 4924
rect 6942 4864 7006 4868
rect 7022 4924 7086 4928
rect 7022 4868 7026 4924
rect 7026 4868 7082 4924
rect 7082 4868 7086 4924
rect 7022 4864 7086 4868
rect 10669 4924 10733 4928
rect 10669 4868 10673 4924
rect 10673 4868 10729 4924
rect 10729 4868 10733 4924
rect 10669 4864 10733 4868
rect 10749 4924 10813 4928
rect 10749 4868 10753 4924
rect 10753 4868 10809 4924
rect 10809 4868 10813 4924
rect 10749 4864 10813 4868
rect 10829 4924 10893 4928
rect 10829 4868 10833 4924
rect 10833 4868 10889 4924
rect 10889 4868 10893 4924
rect 10829 4864 10893 4868
rect 10909 4924 10973 4928
rect 10909 4868 10913 4924
rect 10913 4868 10969 4924
rect 10969 4868 10973 4924
rect 10909 4864 10973 4868
rect 14556 4924 14620 4928
rect 14556 4868 14560 4924
rect 14560 4868 14616 4924
rect 14616 4868 14620 4924
rect 14556 4864 14620 4868
rect 14636 4924 14700 4928
rect 14636 4868 14640 4924
rect 14640 4868 14696 4924
rect 14696 4868 14700 4924
rect 14636 4864 14700 4868
rect 14716 4924 14780 4928
rect 14716 4868 14720 4924
rect 14720 4868 14776 4924
rect 14776 4868 14780 4924
rect 14716 4864 14780 4868
rect 14796 4924 14860 4928
rect 14796 4868 14800 4924
rect 14800 4868 14856 4924
rect 14856 4868 14860 4924
rect 14796 4864 14860 4868
rect 4838 4380 4902 4384
rect 4838 4324 4842 4380
rect 4842 4324 4898 4380
rect 4898 4324 4902 4380
rect 4838 4320 4902 4324
rect 4918 4380 4982 4384
rect 4918 4324 4922 4380
rect 4922 4324 4978 4380
rect 4978 4324 4982 4380
rect 4918 4320 4982 4324
rect 4998 4380 5062 4384
rect 4998 4324 5002 4380
rect 5002 4324 5058 4380
rect 5058 4324 5062 4380
rect 4998 4320 5062 4324
rect 5078 4380 5142 4384
rect 5078 4324 5082 4380
rect 5082 4324 5138 4380
rect 5138 4324 5142 4380
rect 5078 4320 5142 4324
rect 8725 4380 8789 4384
rect 8725 4324 8729 4380
rect 8729 4324 8785 4380
rect 8785 4324 8789 4380
rect 8725 4320 8789 4324
rect 8805 4380 8869 4384
rect 8805 4324 8809 4380
rect 8809 4324 8865 4380
rect 8865 4324 8869 4380
rect 8805 4320 8869 4324
rect 8885 4380 8949 4384
rect 8885 4324 8889 4380
rect 8889 4324 8945 4380
rect 8945 4324 8949 4380
rect 8885 4320 8949 4324
rect 8965 4380 9029 4384
rect 8965 4324 8969 4380
rect 8969 4324 9025 4380
rect 9025 4324 9029 4380
rect 8965 4320 9029 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 16499 4380 16563 4384
rect 16499 4324 16503 4380
rect 16503 4324 16559 4380
rect 16559 4324 16563 4380
rect 16499 4320 16563 4324
rect 16579 4380 16643 4384
rect 16579 4324 16583 4380
rect 16583 4324 16639 4380
rect 16639 4324 16643 4380
rect 16579 4320 16643 4324
rect 16659 4380 16723 4384
rect 16659 4324 16663 4380
rect 16663 4324 16719 4380
rect 16719 4324 16723 4380
rect 16659 4320 16723 4324
rect 16739 4380 16803 4384
rect 16739 4324 16743 4380
rect 16743 4324 16799 4380
rect 16799 4324 16803 4380
rect 16739 4320 16803 4324
rect 2895 3836 2959 3840
rect 2895 3780 2899 3836
rect 2899 3780 2955 3836
rect 2955 3780 2959 3836
rect 2895 3776 2959 3780
rect 2975 3836 3039 3840
rect 2975 3780 2979 3836
rect 2979 3780 3035 3836
rect 3035 3780 3039 3836
rect 2975 3776 3039 3780
rect 3055 3836 3119 3840
rect 3055 3780 3059 3836
rect 3059 3780 3115 3836
rect 3115 3780 3119 3836
rect 3055 3776 3119 3780
rect 3135 3836 3199 3840
rect 3135 3780 3139 3836
rect 3139 3780 3195 3836
rect 3195 3780 3199 3836
rect 3135 3776 3199 3780
rect 6782 3836 6846 3840
rect 6782 3780 6786 3836
rect 6786 3780 6842 3836
rect 6842 3780 6846 3836
rect 6782 3776 6846 3780
rect 6862 3836 6926 3840
rect 6862 3780 6866 3836
rect 6866 3780 6922 3836
rect 6922 3780 6926 3836
rect 6862 3776 6926 3780
rect 6942 3836 7006 3840
rect 6942 3780 6946 3836
rect 6946 3780 7002 3836
rect 7002 3780 7006 3836
rect 6942 3776 7006 3780
rect 7022 3836 7086 3840
rect 7022 3780 7026 3836
rect 7026 3780 7082 3836
rect 7082 3780 7086 3836
rect 7022 3776 7086 3780
rect 10669 3836 10733 3840
rect 10669 3780 10673 3836
rect 10673 3780 10729 3836
rect 10729 3780 10733 3836
rect 10669 3776 10733 3780
rect 10749 3836 10813 3840
rect 10749 3780 10753 3836
rect 10753 3780 10809 3836
rect 10809 3780 10813 3836
rect 10749 3776 10813 3780
rect 10829 3836 10893 3840
rect 10829 3780 10833 3836
rect 10833 3780 10889 3836
rect 10889 3780 10893 3836
rect 10829 3776 10893 3780
rect 10909 3836 10973 3840
rect 10909 3780 10913 3836
rect 10913 3780 10969 3836
rect 10969 3780 10973 3836
rect 10909 3776 10973 3780
rect 14556 3836 14620 3840
rect 14556 3780 14560 3836
rect 14560 3780 14616 3836
rect 14616 3780 14620 3836
rect 14556 3776 14620 3780
rect 14636 3836 14700 3840
rect 14636 3780 14640 3836
rect 14640 3780 14696 3836
rect 14696 3780 14700 3836
rect 14636 3776 14700 3780
rect 14716 3836 14780 3840
rect 14716 3780 14720 3836
rect 14720 3780 14776 3836
rect 14776 3780 14780 3836
rect 14716 3776 14780 3780
rect 14796 3836 14860 3840
rect 14796 3780 14800 3836
rect 14800 3780 14856 3836
rect 14856 3780 14860 3836
rect 14796 3776 14860 3780
rect 4838 3292 4902 3296
rect 4838 3236 4842 3292
rect 4842 3236 4898 3292
rect 4898 3236 4902 3292
rect 4838 3232 4902 3236
rect 4918 3292 4982 3296
rect 4918 3236 4922 3292
rect 4922 3236 4978 3292
rect 4978 3236 4982 3292
rect 4918 3232 4982 3236
rect 4998 3292 5062 3296
rect 4998 3236 5002 3292
rect 5002 3236 5058 3292
rect 5058 3236 5062 3292
rect 4998 3232 5062 3236
rect 5078 3292 5142 3296
rect 5078 3236 5082 3292
rect 5082 3236 5138 3292
rect 5138 3236 5142 3292
rect 5078 3232 5142 3236
rect 8725 3292 8789 3296
rect 8725 3236 8729 3292
rect 8729 3236 8785 3292
rect 8785 3236 8789 3292
rect 8725 3232 8789 3236
rect 8805 3292 8869 3296
rect 8805 3236 8809 3292
rect 8809 3236 8865 3292
rect 8865 3236 8869 3292
rect 8805 3232 8869 3236
rect 8885 3292 8949 3296
rect 8885 3236 8889 3292
rect 8889 3236 8945 3292
rect 8945 3236 8949 3292
rect 8885 3232 8949 3236
rect 8965 3292 9029 3296
rect 8965 3236 8969 3292
rect 8969 3236 9025 3292
rect 9025 3236 9029 3292
rect 8965 3232 9029 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 16499 3292 16563 3296
rect 16499 3236 16503 3292
rect 16503 3236 16559 3292
rect 16559 3236 16563 3292
rect 16499 3232 16563 3236
rect 16579 3292 16643 3296
rect 16579 3236 16583 3292
rect 16583 3236 16639 3292
rect 16639 3236 16643 3292
rect 16579 3232 16643 3236
rect 16659 3292 16723 3296
rect 16659 3236 16663 3292
rect 16663 3236 16719 3292
rect 16719 3236 16723 3292
rect 16659 3232 16723 3236
rect 16739 3292 16803 3296
rect 16739 3236 16743 3292
rect 16743 3236 16799 3292
rect 16799 3236 16803 3292
rect 16739 3232 16803 3236
rect 2895 2748 2959 2752
rect 2895 2692 2899 2748
rect 2899 2692 2955 2748
rect 2955 2692 2959 2748
rect 2895 2688 2959 2692
rect 2975 2748 3039 2752
rect 2975 2692 2979 2748
rect 2979 2692 3035 2748
rect 3035 2692 3039 2748
rect 2975 2688 3039 2692
rect 3055 2748 3119 2752
rect 3055 2692 3059 2748
rect 3059 2692 3115 2748
rect 3115 2692 3119 2748
rect 3055 2688 3119 2692
rect 3135 2748 3199 2752
rect 3135 2692 3139 2748
rect 3139 2692 3195 2748
rect 3195 2692 3199 2748
rect 3135 2688 3199 2692
rect 6782 2748 6846 2752
rect 6782 2692 6786 2748
rect 6786 2692 6842 2748
rect 6842 2692 6846 2748
rect 6782 2688 6846 2692
rect 6862 2748 6926 2752
rect 6862 2692 6866 2748
rect 6866 2692 6922 2748
rect 6922 2692 6926 2748
rect 6862 2688 6926 2692
rect 6942 2748 7006 2752
rect 6942 2692 6946 2748
rect 6946 2692 7002 2748
rect 7002 2692 7006 2748
rect 6942 2688 7006 2692
rect 7022 2748 7086 2752
rect 7022 2692 7026 2748
rect 7026 2692 7082 2748
rect 7082 2692 7086 2748
rect 7022 2688 7086 2692
rect 10669 2748 10733 2752
rect 10669 2692 10673 2748
rect 10673 2692 10729 2748
rect 10729 2692 10733 2748
rect 10669 2688 10733 2692
rect 10749 2748 10813 2752
rect 10749 2692 10753 2748
rect 10753 2692 10809 2748
rect 10809 2692 10813 2748
rect 10749 2688 10813 2692
rect 10829 2748 10893 2752
rect 10829 2692 10833 2748
rect 10833 2692 10889 2748
rect 10889 2692 10893 2748
rect 10829 2688 10893 2692
rect 10909 2748 10973 2752
rect 10909 2692 10913 2748
rect 10913 2692 10969 2748
rect 10969 2692 10973 2748
rect 10909 2688 10973 2692
rect 14556 2748 14620 2752
rect 14556 2692 14560 2748
rect 14560 2692 14616 2748
rect 14616 2692 14620 2748
rect 14556 2688 14620 2692
rect 14636 2748 14700 2752
rect 14636 2692 14640 2748
rect 14640 2692 14696 2748
rect 14696 2692 14700 2748
rect 14636 2688 14700 2692
rect 14716 2748 14780 2752
rect 14716 2692 14720 2748
rect 14720 2692 14776 2748
rect 14776 2692 14780 2748
rect 14716 2688 14780 2692
rect 14796 2748 14860 2752
rect 14796 2692 14800 2748
rect 14800 2692 14856 2748
rect 14856 2692 14860 2748
rect 14796 2688 14860 2692
rect 4838 2204 4902 2208
rect 4838 2148 4842 2204
rect 4842 2148 4898 2204
rect 4898 2148 4902 2204
rect 4838 2144 4902 2148
rect 4918 2204 4982 2208
rect 4918 2148 4922 2204
rect 4922 2148 4978 2204
rect 4978 2148 4982 2204
rect 4918 2144 4982 2148
rect 4998 2204 5062 2208
rect 4998 2148 5002 2204
rect 5002 2148 5058 2204
rect 5058 2148 5062 2204
rect 4998 2144 5062 2148
rect 5078 2204 5142 2208
rect 5078 2148 5082 2204
rect 5082 2148 5138 2204
rect 5138 2148 5142 2204
rect 5078 2144 5142 2148
rect 8725 2204 8789 2208
rect 8725 2148 8729 2204
rect 8729 2148 8785 2204
rect 8785 2148 8789 2204
rect 8725 2144 8789 2148
rect 8805 2204 8869 2208
rect 8805 2148 8809 2204
rect 8809 2148 8865 2204
rect 8865 2148 8869 2204
rect 8805 2144 8869 2148
rect 8885 2204 8949 2208
rect 8885 2148 8889 2204
rect 8889 2148 8945 2204
rect 8945 2148 8949 2204
rect 8885 2144 8949 2148
rect 8965 2204 9029 2208
rect 8965 2148 8969 2204
rect 8969 2148 9025 2204
rect 9025 2148 9029 2204
rect 8965 2144 9029 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 16499 2204 16563 2208
rect 16499 2148 16503 2204
rect 16503 2148 16559 2204
rect 16559 2148 16563 2204
rect 16499 2144 16563 2148
rect 16579 2204 16643 2208
rect 16579 2148 16583 2204
rect 16583 2148 16639 2204
rect 16639 2148 16643 2204
rect 16579 2144 16643 2148
rect 16659 2204 16723 2208
rect 16659 2148 16663 2204
rect 16663 2148 16719 2204
rect 16719 2148 16723 2204
rect 16659 2144 16723 2148
rect 16739 2204 16803 2208
rect 16739 2148 16743 2204
rect 16743 2148 16799 2204
rect 16799 2148 16803 2204
rect 16739 2144 16803 2148
<< metal4 >>
rect 2887 16896 3207 17456
rect 2887 16832 2895 16896
rect 2959 16832 2975 16896
rect 3039 16832 3055 16896
rect 3119 16832 3135 16896
rect 3199 16832 3207 16896
rect 2887 15808 3207 16832
rect 2887 15744 2895 15808
rect 2959 15744 2975 15808
rect 3039 15744 3055 15808
rect 3119 15744 3135 15808
rect 3199 15744 3207 15808
rect 2887 14720 3207 15744
rect 2887 14656 2895 14720
rect 2959 14656 2975 14720
rect 3039 14656 3055 14720
rect 3119 14656 3135 14720
rect 3199 14656 3207 14720
rect 2887 13632 3207 14656
rect 2887 13568 2895 13632
rect 2959 13568 2975 13632
rect 3039 13568 3055 13632
rect 3119 13568 3135 13632
rect 3199 13568 3207 13632
rect 2887 12544 3207 13568
rect 2887 12480 2895 12544
rect 2959 12480 2975 12544
rect 3039 12480 3055 12544
rect 3119 12480 3135 12544
rect 3199 12480 3207 12544
rect 2887 11456 3207 12480
rect 2887 11392 2895 11456
rect 2959 11392 2975 11456
rect 3039 11392 3055 11456
rect 3119 11392 3135 11456
rect 3199 11392 3207 11456
rect 2887 10368 3207 11392
rect 2887 10304 2895 10368
rect 2959 10304 2975 10368
rect 3039 10304 3055 10368
rect 3119 10304 3135 10368
rect 3199 10304 3207 10368
rect 2887 9280 3207 10304
rect 2887 9216 2895 9280
rect 2959 9216 2975 9280
rect 3039 9216 3055 9280
rect 3119 9216 3135 9280
rect 3199 9216 3207 9280
rect 2887 8192 3207 9216
rect 2887 8128 2895 8192
rect 2959 8128 2975 8192
rect 3039 8128 3055 8192
rect 3119 8128 3135 8192
rect 3199 8128 3207 8192
rect 2887 7104 3207 8128
rect 2887 7040 2895 7104
rect 2959 7040 2975 7104
rect 3039 7040 3055 7104
rect 3119 7040 3135 7104
rect 3199 7040 3207 7104
rect 2887 6016 3207 7040
rect 2887 5952 2895 6016
rect 2959 5952 2975 6016
rect 3039 5952 3055 6016
rect 3119 5952 3135 6016
rect 3199 5952 3207 6016
rect 2887 4928 3207 5952
rect 2887 4864 2895 4928
rect 2959 4864 2975 4928
rect 3039 4864 3055 4928
rect 3119 4864 3135 4928
rect 3199 4864 3207 4928
rect 2887 3840 3207 4864
rect 2887 3776 2895 3840
rect 2959 3776 2975 3840
rect 3039 3776 3055 3840
rect 3119 3776 3135 3840
rect 3199 3776 3207 3840
rect 2887 2752 3207 3776
rect 2887 2688 2895 2752
rect 2959 2688 2975 2752
rect 3039 2688 3055 2752
rect 3119 2688 3135 2752
rect 3199 2688 3207 2752
rect 2887 2128 3207 2688
rect 4830 17440 5150 17456
rect 4830 17376 4838 17440
rect 4902 17376 4918 17440
rect 4982 17376 4998 17440
rect 5062 17376 5078 17440
rect 5142 17376 5150 17440
rect 4830 16352 5150 17376
rect 4830 16288 4838 16352
rect 4902 16288 4918 16352
rect 4982 16288 4998 16352
rect 5062 16288 5078 16352
rect 5142 16288 5150 16352
rect 4830 15264 5150 16288
rect 4830 15200 4838 15264
rect 4902 15200 4918 15264
rect 4982 15200 4998 15264
rect 5062 15200 5078 15264
rect 5142 15200 5150 15264
rect 4830 14176 5150 15200
rect 4830 14112 4838 14176
rect 4902 14112 4918 14176
rect 4982 14112 4998 14176
rect 5062 14112 5078 14176
rect 5142 14112 5150 14176
rect 4830 13088 5150 14112
rect 4830 13024 4838 13088
rect 4902 13024 4918 13088
rect 4982 13024 4998 13088
rect 5062 13024 5078 13088
rect 5142 13024 5150 13088
rect 4830 12000 5150 13024
rect 4830 11936 4838 12000
rect 4902 11936 4918 12000
rect 4982 11936 4998 12000
rect 5062 11936 5078 12000
rect 5142 11936 5150 12000
rect 4830 10912 5150 11936
rect 4830 10848 4838 10912
rect 4902 10848 4918 10912
rect 4982 10848 4998 10912
rect 5062 10848 5078 10912
rect 5142 10848 5150 10912
rect 4830 9824 5150 10848
rect 4830 9760 4838 9824
rect 4902 9760 4918 9824
rect 4982 9760 4998 9824
rect 5062 9760 5078 9824
rect 5142 9760 5150 9824
rect 4830 8736 5150 9760
rect 4830 8672 4838 8736
rect 4902 8672 4918 8736
rect 4982 8672 4998 8736
rect 5062 8672 5078 8736
rect 5142 8672 5150 8736
rect 4830 7648 5150 8672
rect 4830 7584 4838 7648
rect 4902 7584 4918 7648
rect 4982 7584 4998 7648
rect 5062 7584 5078 7648
rect 5142 7584 5150 7648
rect 4830 6560 5150 7584
rect 4830 6496 4838 6560
rect 4902 6496 4918 6560
rect 4982 6496 4998 6560
rect 5062 6496 5078 6560
rect 5142 6496 5150 6560
rect 4830 5472 5150 6496
rect 4830 5408 4838 5472
rect 4902 5408 4918 5472
rect 4982 5408 4998 5472
rect 5062 5408 5078 5472
rect 5142 5408 5150 5472
rect 4830 4384 5150 5408
rect 4830 4320 4838 4384
rect 4902 4320 4918 4384
rect 4982 4320 4998 4384
rect 5062 4320 5078 4384
rect 5142 4320 5150 4384
rect 4830 3296 5150 4320
rect 4830 3232 4838 3296
rect 4902 3232 4918 3296
rect 4982 3232 4998 3296
rect 5062 3232 5078 3296
rect 5142 3232 5150 3296
rect 4830 2208 5150 3232
rect 4830 2144 4838 2208
rect 4902 2144 4918 2208
rect 4982 2144 4998 2208
rect 5062 2144 5078 2208
rect 5142 2144 5150 2208
rect 4830 2128 5150 2144
rect 6774 16896 7094 17456
rect 6774 16832 6782 16896
rect 6846 16832 6862 16896
rect 6926 16832 6942 16896
rect 7006 16832 7022 16896
rect 7086 16832 7094 16896
rect 6774 15808 7094 16832
rect 6774 15744 6782 15808
rect 6846 15744 6862 15808
rect 6926 15744 6942 15808
rect 7006 15744 7022 15808
rect 7086 15744 7094 15808
rect 6774 14720 7094 15744
rect 6774 14656 6782 14720
rect 6846 14656 6862 14720
rect 6926 14656 6942 14720
rect 7006 14656 7022 14720
rect 7086 14656 7094 14720
rect 6774 13632 7094 14656
rect 6774 13568 6782 13632
rect 6846 13568 6862 13632
rect 6926 13568 6942 13632
rect 7006 13568 7022 13632
rect 7086 13568 7094 13632
rect 6774 12544 7094 13568
rect 6774 12480 6782 12544
rect 6846 12480 6862 12544
rect 6926 12480 6942 12544
rect 7006 12480 7022 12544
rect 7086 12480 7094 12544
rect 6774 11456 7094 12480
rect 6774 11392 6782 11456
rect 6846 11392 6862 11456
rect 6926 11392 6942 11456
rect 7006 11392 7022 11456
rect 7086 11392 7094 11456
rect 6774 10368 7094 11392
rect 6774 10304 6782 10368
rect 6846 10304 6862 10368
rect 6926 10304 6942 10368
rect 7006 10304 7022 10368
rect 7086 10304 7094 10368
rect 6774 9280 7094 10304
rect 6774 9216 6782 9280
rect 6846 9216 6862 9280
rect 6926 9216 6942 9280
rect 7006 9216 7022 9280
rect 7086 9216 7094 9280
rect 6774 8192 7094 9216
rect 6774 8128 6782 8192
rect 6846 8128 6862 8192
rect 6926 8128 6942 8192
rect 7006 8128 7022 8192
rect 7086 8128 7094 8192
rect 6774 7104 7094 8128
rect 6774 7040 6782 7104
rect 6846 7040 6862 7104
rect 6926 7040 6942 7104
rect 7006 7040 7022 7104
rect 7086 7040 7094 7104
rect 6774 6016 7094 7040
rect 6774 5952 6782 6016
rect 6846 5952 6862 6016
rect 6926 5952 6942 6016
rect 7006 5952 7022 6016
rect 7086 5952 7094 6016
rect 6774 4928 7094 5952
rect 6774 4864 6782 4928
rect 6846 4864 6862 4928
rect 6926 4864 6942 4928
rect 7006 4864 7022 4928
rect 7086 4864 7094 4928
rect 6774 3840 7094 4864
rect 6774 3776 6782 3840
rect 6846 3776 6862 3840
rect 6926 3776 6942 3840
rect 7006 3776 7022 3840
rect 7086 3776 7094 3840
rect 6774 2752 7094 3776
rect 6774 2688 6782 2752
rect 6846 2688 6862 2752
rect 6926 2688 6942 2752
rect 7006 2688 7022 2752
rect 7086 2688 7094 2752
rect 6774 2128 7094 2688
rect 8717 17440 9037 17456
rect 8717 17376 8725 17440
rect 8789 17376 8805 17440
rect 8869 17376 8885 17440
rect 8949 17376 8965 17440
rect 9029 17376 9037 17440
rect 8717 16352 9037 17376
rect 8717 16288 8725 16352
rect 8789 16288 8805 16352
rect 8869 16288 8885 16352
rect 8949 16288 8965 16352
rect 9029 16288 9037 16352
rect 8717 15264 9037 16288
rect 8717 15200 8725 15264
rect 8789 15200 8805 15264
rect 8869 15200 8885 15264
rect 8949 15200 8965 15264
rect 9029 15200 9037 15264
rect 8717 14176 9037 15200
rect 8717 14112 8725 14176
rect 8789 14112 8805 14176
rect 8869 14112 8885 14176
rect 8949 14112 8965 14176
rect 9029 14112 9037 14176
rect 8717 13088 9037 14112
rect 8717 13024 8725 13088
rect 8789 13024 8805 13088
rect 8869 13024 8885 13088
rect 8949 13024 8965 13088
rect 9029 13024 9037 13088
rect 8717 12000 9037 13024
rect 8717 11936 8725 12000
rect 8789 11936 8805 12000
rect 8869 11936 8885 12000
rect 8949 11936 8965 12000
rect 9029 11936 9037 12000
rect 8717 10912 9037 11936
rect 8717 10848 8725 10912
rect 8789 10848 8805 10912
rect 8869 10848 8885 10912
rect 8949 10848 8965 10912
rect 9029 10848 9037 10912
rect 8717 9824 9037 10848
rect 8717 9760 8725 9824
rect 8789 9760 8805 9824
rect 8869 9760 8885 9824
rect 8949 9760 8965 9824
rect 9029 9760 9037 9824
rect 8717 8736 9037 9760
rect 8717 8672 8725 8736
rect 8789 8672 8805 8736
rect 8869 8672 8885 8736
rect 8949 8672 8965 8736
rect 9029 8672 9037 8736
rect 8717 7648 9037 8672
rect 8717 7584 8725 7648
rect 8789 7584 8805 7648
rect 8869 7584 8885 7648
rect 8949 7584 8965 7648
rect 9029 7584 9037 7648
rect 8717 6560 9037 7584
rect 8717 6496 8725 6560
rect 8789 6496 8805 6560
rect 8869 6496 8885 6560
rect 8949 6496 8965 6560
rect 9029 6496 9037 6560
rect 8717 5472 9037 6496
rect 8717 5408 8725 5472
rect 8789 5408 8805 5472
rect 8869 5408 8885 5472
rect 8949 5408 8965 5472
rect 9029 5408 9037 5472
rect 8717 4384 9037 5408
rect 8717 4320 8725 4384
rect 8789 4320 8805 4384
rect 8869 4320 8885 4384
rect 8949 4320 8965 4384
rect 9029 4320 9037 4384
rect 8717 3296 9037 4320
rect 8717 3232 8725 3296
rect 8789 3232 8805 3296
rect 8869 3232 8885 3296
rect 8949 3232 8965 3296
rect 9029 3232 9037 3296
rect 8717 2208 9037 3232
rect 8717 2144 8725 2208
rect 8789 2144 8805 2208
rect 8869 2144 8885 2208
rect 8949 2144 8965 2208
rect 9029 2144 9037 2208
rect 8717 2128 9037 2144
rect 10661 16896 10981 17456
rect 10661 16832 10669 16896
rect 10733 16832 10749 16896
rect 10813 16832 10829 16896
rect 10893 16832 10909 16896
rect 10973 16832 10981 16896
rect 10661 15808 10981 16832
rect 10661 15744 10669 15808
rect 10733 15744 10749 15808
rect 10813 15744 10829 15808
rect 10893 15744 10909 15808
rect 10973 15744 10981 15808
rect 10661 14720 10981 15744
rect 10661 14656 10669 14720
rect 10733 14656 10749 14720
rect 10813 14656 10829 14720
rect 10893 14656 10909 14720
rect 10973 14656 10981 14720
rect 10661 13632 10981 14656
rect 10661 13568 10669 13632
rect 10733 13568 10749 13632
rect 10813 13568 10829 13632
rect 10893 13568 10909 13632
rect 10973 13568 10981 13632
rect 10661 12544 10981 13568
rect 10661 12480 10669 12544
rect 10733 12480 10749 12544
rect 10813 12480 10829 12544
rect 10893 12480 10909 12544
rect 10973 12480 10981 12544
rect 10661 11456 10981 12480
rect 10661 11392 10669 11456
rect 10733 11392 10749 11456
rect 10813 11392 10829 11456
rect 10893 11392 10909 11456
rect 10973 11392 10981 11456
rect 10661 10368 10981 11392
rect 10661 10304 10669 10368
rect 10733 10304 10749 10368
rect 10813 10304 10829 10368
rect 10893 10304 10909 10368
rect 10973 10304 10981 10368
rect 10661 9280 10981 10304
rect 10661 9216 10669 9280
rect 10733 9216 10749 9280
rect 10813 9216 10829 9280
rect 10893 9216 10909 9280
rect 10973 9216 10981 9280
rect 10661 8192 10981 9216
rect 10661 8128 10669 8192
rect 10733 8128 10749 8192
rect 10813 8128 10829 8192
rect 10893 8128 10909 8192
rect 10973 8128 10981 8192
rect 10661 7104 10981 8128
rect 10661 7040 10669 7104
rect 10733 7040 10749 7104
rect 10813 7040 10829 7104
rect 10893 7040 10909 7104
rect 10973 7040 10981 7104
rect 10661 6016 10981 7040
rect 10661 5952 10669 6016
rect 10733 5952 10749 6016
rect 10813 5952 10829 6016
rect 10893 5952 10909 6016
rect 10973 5952 10981 6016
rect 10661 4928 10981 5952
rect 10661 4864 10669 4928
rect 10733 4864 10749 4928
rect 10813 4864 10829 4928
rect 10893 4864 10909 4928
rect 10973 4864 10981 4928
rect 10661 3840 10981 4864
rect 10661 3776 10669 3840
rect 10733 3776 10749 3840
rect 10813 3776 10829 3840
rect 10893 3776 10909 3840
rect 10973 3776 10981 3840
rect 10661 2752 10981 3776
rect 10661 2688 10669 2752
rect 10733 2688 10749 2752
rect 10813 2688 10829 2752
rect 10893 2688 10909 2752
rect 10973 2688 10981 2752
rect 10661 2128 10981 2688
rect 12604 17440 12924 17456
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13088 12924 14112
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12604 8736 12924 9760
rect 12604 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3296 12924 4320
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 14548 16896 14868 17456
rect 14548 16832 14556 16896
rect 14620 16832 14636 16896
rect 14700 16832 14716 16896
rect 14780 16832 14796 16896
rect 14860 16832 14868 16896
rect 14548 15808 14868 16832
rect 14548 15744 14556 15808
rect 14620 15744 14636 15808
rect 14700 15744 14716 15808
rect 14780 15744 14796 15808
rect 14860 15744 14868 15808
rect 14548 14720 14868 15744
rect 14548 14656 14556 14720
rect 14620 14656 14636 14720
rect 14700 14656 14716 14720
rect 14780 14656 14796 14720
rect 14860 14656 14868 14720
rect 14548 13632 14868 14656
rect 14548 13568 14556 13632
rect 14620 13568 14636 13632
rect 14700 13568 14716 13632
rect 14780 13568 14796 13632
rect 14860 13568 14868 13632
rect 14548 12544 14868 13568
rect 14548 12480 14556 12544
rect 14620 12480 14636 12544
rect 14700 12480 14716 12544
rect 14780 12480 14796 12544
rect 14860 12480 14868 12544
rect 14548 11456 14868 12480
rect 14548 11392 14556 11456
rect 14620 11392 14636 11456
rect 14700 11392 14716 11456
rect 14780 11392 14796 11456
rect 14860 11392 14868 11456
rect 14548 10368 14868 11392
rect 14548 10304 14556 10368
rect 14620 10304 14636 10368
rect 14700 10304 14716 10368
rect 14780 10304 14796 10368
rect 14860 10304 14868 10368
rect 14548 9280 14868 10304
rect 14548 9216 14556 9280
rect 14620 9216 14636 9280
rect 14700 9216 14716 9280
rect 14780 9216 14796 9280
rect 14860 9216 14868 9280
rect 14548 8192 14868 9216
rect 14548 8128 14556 8192
rect 14620 8128 14636 8192
rect 14700 8128 14716 8192
rect 14780 8128 14796 8192
rect 14860 8128 14868 8192
rect 14548 7104 14868 8128
rect 14548 7040 14556 7104
rect 14620 7040 14636 7104
rect 14700 7040 14716 7104
rect 14780 7040 14796 7104
rect 14860 7040 14868 7104
rect 14548 6016 14868 7040
rect 14548 5952 14556 6016
rect 14620 5952 14636 6016
rect 14700 5952 14716 6016
rect 14780 5952 14796 6016
rect 14860 5952 14868 6016
rect 14548 4928 14868 5952
rect 14548 4864 14556 4928
rect 14620 4864 14636 4928
rect 14700 4864 14716 4928
rect 14780 4864 14796 4928
rect 14860 4864 14868 4928
rect 14548 3840 14868 4864
rect 14548 3776 14556 3840
rect 14620 3776 14636 3840
rect 14700 3776 14716 3840
rect 14780 3776 14796 3840
rect 14860 3776 14868 3840
rect 14548 2752 14868 3776
rect 14548 2688 14556 2752
rect 14620 2688 14636 2752
rect 14700 2688 14716 2752
rect 14780 2688 14796 2752
rect 14860 2688 14868 2752
rect 14548 2128 14868 2688
rect 16491 17440 16811 17456
rect 16491 17376 16499 17440
rect 16563 17376 16579 17440
rect 16643 17376 16659 17440
rect 16723 17376 16739 17440
rect 16803 17376 16811 17440
rect 16491 16352 16811 17376
rect 16491 16288 16499 16352
rect 16563 16288 16579 16352
rect 16643 16288 16659 16352
rect 16723 16288 16739 16352
rect 16803 16288 16811 16352
rect 16491 15264 16811 16288
rect 16491 15200 16499 15264
rect 16563 15200 16579 15264
rect 16643 15200 16659 15264
rect 16723 15200 16739 15264
rect 16803 15200 16811 15264
rect 16491 14176 16811 15200
rect 16491 14112 16499 14176
rect 16563 14112 16579 14176
rect 16643 14112 16659 14176
rect 16723 14112 16739 14176
rect 16803 14112 16811 14176
rect 16491 13088 16811 14112
rect 16491 13024 16499 13088
rect 16563 13024 16579 13088
rect 16643 13024 16659 13088
rect 16723 13024 16739 13088
rect 16803 13024 16811 13088
rect 16491 12000 16811 13024
rect 16491 11936 16499 12000
rect 16563 11936 16579 12000
rect 16643 11936 16659 12000
rect 16723 11936 16739 12000
rect 16803 11936 16811 12000
rect 16491 10912 16811 11936
rect 16491 10848 16499 10912
rect 16563 10848 16579 10912
rect 16643 10848 16659 10912
rect 16723 10848 16739 10912
rect 16803 10848 16811 10912
rect 16491 9824 16811 10848
rect 16491 9760 16499 9824
rect 16563 9760 16579 9824
rect 16643 9760 16659 9824
rect 16723 9760 16739 9824
rect 16803 9760 16811 9824
rect 16491 8736 16811 9760
rect 16491 8672 16499 8736
rect 16563 8672 16579 8736
rect 16643 8672 16659 8736
rect 16723 8672 16739 8736
rect 16803 8672 16811 8736
rect 16491 7648 16811 8672
rect 16491 7584 16499 7648
rect 16563 7584 16579 7648
rect 16643 7584 16659 7648
rect 16723 7584 16739 7648
rect 16803 7584 16811 7648
rect 16491 6560 16811 7584
rect 16491 6496 16499 6560
rect 16563 6496 16579 6560
rect 16643 6496 16659 6560
rect 16723 6496 16739 6560
rect 16803 6496 16811 6560
rect 16491 5472 16811 6496
rect 16491 5408 16499 5472
rect 16563 5408 16579 5472
rect 16643 5408 16659 5472
rect 16723 5408 16739 5472
rect 16803 5408 16811 5472
rect 16491 4384 16811 5408
rect 16491 4320 16499 4384
rect 16563 4320 16579 4384
rect 16643 4320 16659 4384
rect 16723 4320 16739 4384
rect 16803 4320 16811 4384
rect 16491 3296 16811 4320
rect 16491 3232 16499 3296
rect 16563 3232 16579 3296
rect 16643 3232 16659 3296
rect 16723 3232 16739 3296
rect 16803 3232 16811 3296
rect 16491 2208 16811 3232
rect 16491 2144 16499 2208
rect 16563 2144 16579 2208
rect 16643 2144 16659 2208
rect 16723 2144 16739 2208
rect 16803 2144 16811 2208
rect 16491 2128 16811 2144
use sky130_fd_sc_hd__clkbuf_4  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _170_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1688980957
transform 1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _172_
timestamp 1688980957
transform 1 0 5244 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1688980957
transform 1 0 3864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _174_
timestamp 1688980957
transform 1 0 5244 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1688980957
transform 1 0 4784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _176_
timestamp 1688980957
transform 1 0 6992 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _177_
timestamp 1688980957
transform 1 0 6440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _178_
timestamp 1688980957
transform 1 0 4692 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1688980957
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _180_
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _182_
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1688980957
transform 1 0 3220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _185_
timestamp 1688980957
transform 1 0 6164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _186_
timestamp 1688980957
transform 1 0 9016 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _187_
timestamp 1688980957
transform 1 0 9108 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1688980957
transform 1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _189_
timestamp 1688980957
transform 1 0 11960 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _191_
timestamp 1688980957
transform 1 0 10304 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1688980957
transform 1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1688980957
transform 1 0 12696 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1688980957
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1688980957
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _197_
timestamp 1688980957
transform 1 0 14260 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _199_
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp 1688980957
transform 1 0 12604 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1688980957
transform 1 0 12696 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp 1688980957
transform 1 0 14168 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1688980957
transform 1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 1688980957
transform 1 0 14352 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1688980957
transform 1 0 15088 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _207_
timestamp 1688980957
transform 1 0 8832 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1688980957
transform 1 0 14628 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 1688980957
transform 1 0 13340 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1688980957
transform 1 0 12788 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1688980957
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1688980957
transform 1 0 9936 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1688980957
transform 1 0 9752 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1688980957
transform 1 0 7268 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 1688980957
transform 1 0 5428 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1688980957
transform 1 0 5704 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1688980957
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1688980957
transform 1 0 5244 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1688980957
transform 1 0 6440 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _226_
timestamp 1688980957
transform 1 0 7360 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1688980957
transform 1 0 4324 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1688980957
transform 1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1688980957
transform 1 0 2668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1688980957
transform 1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4600 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4600 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _234_
timestamp 1688980957
transform 1 0 5152 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _235_
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1688980957
transform 1 0 1840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7912 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8372 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_4  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _243_
timestamp 1688980957
transform 1 0 6992 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1688980957
transform 1 0 6808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _245_
timestamp 1688980957
transform 1 0 3864 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _246_
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1688980957
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _248_
timestamp 1688980957
transform 1 0 2668 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _249_
timestamp 1688980957
transform 1 0 1840 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1688980957
transform 1 0 1564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _251_
timestamp 1688980957
transform 1 0 8740 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _252_
timestamp 1688980957
transform 1 0 7912 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1688980957
transform 1 0 6992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _254_
timestamp 1688980957
transform 1 0 5060 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _255_
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1688980957
transform 1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _257_
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _258_
timestamp 1688980957
transform 1 0 5336 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1688980957
transform 1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _260_
timestamp 1688980957
transform 1 0 2760 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _261_
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1688980957
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _263_
timestamp 1688980957
transform 1 0 2024 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _264_
timestamp 1688980957
transform 1 0 1840 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp 1688980957
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10396 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _270_
timestamp 1688980957
transform 1 0 11500 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _273_
timestamp 1688980957
transform 1 0 11684 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _274_
timestamp 1688980957
transform 1 0 11592 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _275_
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _276_
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _277_
timestamp 1688980957
transform 1 0 10488 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _278_
timestamp 1688980957
transform 1 0 9200 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _279_
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1688980957
transform 1 0 7820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _282_
timestamp 1688980957
transform 1 0 8004 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _283_
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1688980957
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9292 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _286_
timestamp 1688980957
transform 1 0 3404 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_4  _287_
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _288_
timestamp 1688980957
transform 1 0 2576 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 1688980957
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _290_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _291_
timestamp 1688980957
transform 1 0 2852 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1688980957
transform 1 0 2392 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _293_
timestamp 1688980957
transform 1 0 3220 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _294_
timestamp 1688980957
transform 1 0 3404 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp 1688980957
transform 1 0 2944 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _296_
timestamp 1688980957
transform 1 0 8924 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1688980957
transform 1 0 7820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _299_
timestamp 1688980957
transform 1 0 9016 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _300_
timestamp 1688980957
transform 1 0 8924 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp 1688980957
transform 1 0 9752 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _302_
timestamp 1688980957
transform 1 0 4784 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp 1688980957
transform 1 0 4232 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1688980957
transform 1 0 3864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _305_
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 1688980957
transform 1 0 6072 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1688980957
transform 1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _308_
timestamp 1688980957
transform 1 0 7084 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _309_
timestamp 1688980957
transform 1 0 6992 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1688980957
transform 1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _312_
timestamp 1688980957
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10396 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _314_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _315_
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _316_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _317_
timestamp 1688980957
transform 1 0 11776 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _318_
timestamp 1688980957
transform 1 0 12328 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _319_
timestamp 1688980957
transform 1 0 11960 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _320_
timestamp 1688980957
transform 1 0 11592 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _321_
timestamp 1688980957
transform 1 0 11868 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _322_
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _323_
timestamp 1688980957
transform 1 0 15364 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1688980957
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _326_
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1688980957
transform 1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9568 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1688980957
transform 1 0 9108 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1688980957
transform 1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _331_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1688980957
transform 1 0 4416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1688980957
transform 1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1688980957
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1688980957
transform 1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1688980957
transform 1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1688980957
transform 1 0 3864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1688980957
transform 1 0 6716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _342_
timestamp 1688980957
transform 1 0 10672 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1688980957
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1688980957
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1688980957
transform 1 0 15548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1688980957
transform 1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1688980957
transform 1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1688980957
transform 1 0 13616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1688980957
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1688980957
transform 1 0 15272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _353_
timestamp 1688980957
transform 1 0 10212 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1688980957
transform 1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1688980957
transform 1 0 12144 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1688980957
transform 1 0 10580 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1688980957
transform 1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1688980957
transform 1 0 6808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1688980957
transform 1 0 6164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1688980957
transform 1 0 6900 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1688980957
transform 1 0 8280 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1688980957
transform 1 0 7452 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1688980957
transform 1 0 3864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1688980957
transform 1 0 2300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _366_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _367_
timestamp 1688980957
transform 1 0 2392 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _369_
timestamp 1688980957
transform 1 0 6440 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _372_
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _373_
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _374_
timestamp 1688980957
transform 1 0 11960 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _375_
timestamp 1688980957
transform 1 0 12328 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _376_
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _377_
timestamp 1688980957
transform 1 0 11960 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _378_
timestamp 1688980957
transform 1 0 9752 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _379_
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1688980957
transform 1 0 8648 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _381_
timestamp 1688980957
transform 1 0 8464 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1688980957
transform 1 0 1656 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _387_
timestamp 1688980957
transform 1 0 9016 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1688980957
transform 1 0 3772 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1688980957
transform 1 0 4600 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1688980957
transform 1 0 6532 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1688980957
transform 1 0 10764 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1688980957
transform 1 0 10764 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1688980957
transform 1 0 11776 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1688980957
transform 1 0 12880 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1688980957
transform 1 0 12512 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _398_
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _401_
timestamp 1688980957
transform 1 0 9200 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _402_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1688980957
transform 1 0 2576 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _404_
timestamp 1688980957
transform 1 0 3128 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _405_
timestamp 1688980957
transform 1 0 4232 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _406_
timestamp 1688980957
transform 1 0 6716 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _407_
timestamp 1688980957
transform 1 0 5520 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _408_
timestamp 1688980957
transform 1 0 3404 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _409_
timestamp 1688980957
transform 1 0 2668 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _410_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _411_
timestamp 1688980957
transform 1 0 6992 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _412_
timestamp 1688980957
transform 1 0 10120 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _413_
timestamp 1688980957
transform 1 0 9568 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _414_
timestamp 1688980957
transform 1 0 11868 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _415_
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _416_
timestamp 1688980957
transform 1 0 14168 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _417_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _418_
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _419_
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _420_
timestamp 1688980957
transform 1 0 14444 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _421_
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _422_
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _423_
timestamp 1688980957
transform 1 0 12880 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _424_
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _425_
timestamp 1688980957
transform 1 0 9568 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _426_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _427_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _428_
timestamp 1688980957
transform 1 0 4416 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _429_
timestamp 1688980957
transform 1 0 5152 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _430_
timestamp 1688980957
transform 1 0 6992 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _431_
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _432_
timestamp 1688980957
transform 1 0 2852 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _433_
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1688980957
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1688980957
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1688980957
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1688980957
transform 1 0 6440 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 1688980957
transform 1 0 8188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1688980957
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_67
timestamp 1688980957
transform 1 0 7268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_93 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103
timestamp 1688980957
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_127
timestamp 1688980957
transform 1 0 12788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_161
timestamp 1688980957
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_11
timestamp 1688980957
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_35
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_52
timestamp 1688980957
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_88
timestamp 1688980957
transform 1 0 9200 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_117
timestamp 1688980957
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_134
timestamp 1688980957
transform 1 0 13432 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_146
timestamp 1688980957
transform 1 0 14536 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_158
timestamp 1688980957
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_21
timestamp 1688980957
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_38
timestamp 1688980957
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_42
timestamp 1688980957
transform 1 0 4968 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_48
timestamp 1688980957
transform 1 0 5520 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_60
timestamp 1688980957
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_73
timestamp 1688980957
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 1688980957
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_149
timestamp 1688980957
transform 1 0 14812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_161
timestamp 1688980957
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_7
timestamp 1688980957
transform 1 0 1748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_19
timestamp 1688980957
transform 1 0 2852 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_89
timestamp 1688980957
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_116
timestamp 1688980957
transform 1 0 11776 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_135
timestamp 1688980957
transform 1 0 13524 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_160
timestamp 1688980957
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp 1688980957
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_32
timestamp 1688980957
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_38
timestamp 1688980957
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_74
timestamp 1688980957
transform 1 0 7912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1688980957
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_95
timestamp 1688980957
transform 1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_101
timestamp 1688980957
transform 1 0 10396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_113
timestamp 1688980957
transform 1 0 11500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_125
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_150
timestamp 1688980957
transform 1 0 14904 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_162
timestamp 1688980957
transform 1 0 16008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_37
timestamp 1688980957
transform 1 0 4508 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_48
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_76
timestamp 1688980957
transform 1 0 8096 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_98
timestamp 1688980957
transform 1 0 10120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_141
timestamp 1688980957
transform 1 0 14076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_165
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 1688980957
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_33
timestamp 1688980957
transform 1 0 4140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_39
timestamp 1688980957
transform 1 0 4692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_43
timestamp 1688980957
transform 1 0 5060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_48
timestamp 1688980957
transform 1 0 5520 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_54
timestamp 1688980957
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_58
timestamp 1688980957
transform 1 0 6440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_96
timestamp 1688980957
transform 1 0 9936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_130
timestamp 1688980957
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1688980957
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_147
timestamp 1688980957
transform 1 0 14628 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_159
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_26
timestamp 1688980957
transform 1 0 3496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_77
timestamp 1688980957
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_85
timestamp 1688980957
transform 1 0 8924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_97
timestamp 1688980957
transform 1 0 10028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1688980957
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_138
timestamp 1688980957
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_142
timestamp 1688980957
transform 1 0 14168 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_152
timestamp 1688980957
transform 1 0 15088 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_164
timestamp 1688980957
transform 1 0 16192 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_23
timestamp 1688980957
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_33
timestamp 1688980957
transform 1 0 4140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_45
timestamp 1688980957
transform 1 0 5244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_55
timestamp 1688980957
transform 1 0 6164 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_72
timestamp 1688980957
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_94
timestamp 1688980957
transform 1 0 9752 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_161
timestamp 1688980957
transform 1 0 15916 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_19
timestamp 1688980957
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1688980957
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_63
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_73
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_79
timestamp 1688980957
transform 1 0 8372 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_117
timestamp 1688980957
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_134
timestamp 1688980957
transform 1 0 13432 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_139
timestamp 1688980957
transform 1 0 13892 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_143
timestamp 1688980957
transform 1 0 14260 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_154
timestamp 1688980957
transform 1 0 15272 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_19
timestamp 1688980957
transform 1 0 2852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_23
timestamp 1688980957
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_38
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_55
timestamp 1688980957
transform 1 0 6164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_79
timestamp 1688980957
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_100
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_110
timestamp 1688980957
transform 1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_150
timestamp 1688980957
transform 1 0 14904 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_162
timestamp 1688980957
transform 1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_6
timestamp 1688980957
transform 1 0 1656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_36
timestamp 1688980957
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_61
timestamp 1688980957
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_65
timestamp 1688980957
transform 1 0 7084 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_77
timestamp 1688980957
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_96
timestamp 1688980957
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_129
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_153
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_165
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_17
timestamp 1688980957
transform 1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 1688980957
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_33
timestamp 1688980957
transform 1 0 4140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_52
timestamp 1688980957
transform 1 0 5888 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_64
timestamp 1688980957
transform 1 0 6992 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_72
timestamp 1688980957
transform 1 0 7728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_76
timestamp 1688980957
transform 1 0 8096 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_118
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_124
timestamp 1688980957
transform 1 0 12512 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_134
timestamp 1688980957
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_164
timestamp 1688980957
transform 1 0 16192 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_19
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_25
timestamp 1688980957
transform 1 0 3404 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_35
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_62
timestamp 1688980957
transform 1 0 6808 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_66
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_92
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_101
timestamp 1688980957
transform 1 0 10396 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_129
timestamp 1688980957
transform 1 0 12972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_157
timestamp 1688980957
transform 1 0 15548 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_23
timestamp 1688980957
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_55
timestamp 1688980957
transform 1 0 6164 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 1688980957
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1688980957
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_114
timestamp 1688980957
transform 1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_28
timestamp 1688980957
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_38
timestamp 1688980957
transform 1 0 4600 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_45
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_52
timestamp 1688980957
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_61
timestamp 1688980957
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_70
timestamp 1688980957
transform 1 0 7544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_74
timestamp 1688980957
transform 1 0 7912 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_97
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_117
timestamp 1688980957
transform 1 0 11868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_129
timestamp 1688980957
transform 1 0 12972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_141
timestamp 1688980957
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_155
timestamp 1688980957
transform 1 0 15364 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_163
timestamp 1688980957
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_25
timestamp 1688980957
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_34
timestamp 1688980957
transform 1 0 4232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_63
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_73
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_96
timestamp 1688980957
transform 1 0 9936 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_110
timestamp 1688980957
transform 1 0 11224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1688980957
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_161
timestamp 1688980957
transform 1 0 15916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_11
timestamp 1688980957
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_17
timestamp 1688980957
transform 1 0 2668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_29
timestamp 1688980957
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_41
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1688980957
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_75
timestamp 1688980957
transform 1 0 8004 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_87
timestamp 1688980957
transform 1 0 9108 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_91
timestamp 1688980957
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_103
timestamp 1688980957
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_120
timestamp 1688980957
transform 1 0 12144 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_132
timestamp 1688980957
transform 1 0 13248 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_136
timestamp 1688980957
transform 1 0 13616 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_157
timestamp 1688980957
transform 1 0 15548 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_165
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_23
timestamp 1688980957
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_33
timestamp 1688980957
transform 1 0 4140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1688980957
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_45
timestamp 1688980957
transform 1 0 5244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_49
timestamp 1688980957
transform 1 0 5612 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_61
timestamp 1688980957
transform 1 0 6716 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_76
timestamp 1688980957
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_144
timestamp 1688980957
transform 1 0 14352 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_156
timestamp 1688980957
transform 1 0 15456 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_164
timestamp 1688980957
transform 1 0 16192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_9
timestamp 1688980957
transform 1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_117
timestamp 1688980957
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_147
timestamp 1688980957
transform 1 0 14628 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_159
timestamp 1688980957
transform 1 0 15732 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_165
timestamp 1688980957
transform 1 0 16284 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1688980957
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_37
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_45
timestamp 1688980957
transform 1 0 5244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_57
timestamp 1688980957
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_69
timestamp 1688980957
transform 1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_73
timestamp 1688980957
transform 1 0 7820 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_129
timestamp 1688980957
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1688980957
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_161
timestamp 1688980957
transform 1 0 15916 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_7
timestamp 1688980957
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_11
timestamp 1688980957
transform 1 0 2116 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_21
timestamp 1688980957
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_34
timestamp 1688980957
transform 1 0 4232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_90
timestamp 1688980957
transform 1 0 9384 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_123
timestamp 1688980957
transform 1 0 12420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_127
timestamp 1688980957
transform 1 0 12788 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_150
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_18
timestamp 1688980957
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_48
timestamp 1688980957
transform 1 0 5520 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_72
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_76
timestamp 1688980957
transform 1 0 8096 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_106
timestamp 1688980957
transform 1 0 10856 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_114
timestamp 1688980957
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_132
timestamp 1688980957
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_150
timestamp 1688980957
transform 1 0 14904 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_162
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_19
timestamp 1688980957
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_31
timestamp 1688980957
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_43
timestamp 1688980957
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_65
timestamp 1688980957
transform 1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_89
timestamp 1688980957
transform 1 0 9292 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_122
timestamp 1688980957
transform 1 0 12328 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_148
timestamp 1688980957
transform 1 0 14720 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_160
timestamp 1688980957
transform 1 0 15824 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_37
timestamp 1688980957
transform 1 0 4508 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_48
timestamp 1688980957
transform 1 0 5520 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_54
timestamp 1688980957
transform 1 0 6072 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_58
timestamp 1688980957
transform 1 0 6440 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_70
timestamp 1688980957
transform 1 0 7544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1688980957
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_91
timestamp 1688980957
transform 1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_95
timestamp 1688980957
transform 1 0 9844 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_107
timestamp 1688980957
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_119
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_123
timestamp 1688980957
transform 1 0 12420 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_130
timestamp 1688980957
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1688980957
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_144
timestamp 1688980957
transform 1 0 14352 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_156
timestamp 1688980957
transform 1 0 15456 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_164
timestamp 1688980957
transform 1 0 16192 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_14
timestamp 1688980957
transform 1 0 2392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_30
timestamp 1688980957
transform 1 0 3864 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_61
timestamp 1688980957
transform 1 0 6716 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_66
timestamp 1688980957
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_72
timestamp 1688980957
transform 1 0 7728 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_97
timestamp 1688980957
transform 1 0 10028 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_142
timestamp 1688980957
transform 1 0 14168 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_154
timestamp 1688980957
transform 1 0 15272 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_22
timestamp 1688980957
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_33
timestamp 1688980957
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_43
timestamp 1688980957
transform 1 0 5060 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_102
timestamp 1688980957
transform 1 0 10488 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_114
timestamp 1688980957
transform 1 0 11592 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_126
timestamp 1688980957
transform 1 0 12696 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1688980957
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_9
timestamp 1688980957
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_21
timestamp 1688980957
transform 1 0 3036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 1688980957
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_77
timestamp 1688980957
transform 1 0 8188 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_83
timestamp 1688980957
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_94
timestamp 1688980957
transform 1 0 9752 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_106
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_119
timestamp 1688980957
transform 1 0 12052 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_131
timestamp 1688980957
transform 1 0 13156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_139
timestamp 1688980957
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_141
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_153
timestamp 1688980957
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 16100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1688980957
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1688980957
transform 1 0 15824 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1688980957
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1688980957
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1688980957
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1688980957
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1688980957
transform 1 0 7820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 15548 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1688980957
transform -1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1688980957
transform -1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1688980957
transform -1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1688980957
transform -1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1688980957
transform -1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1688980957
transform -1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1688980957
transform -1 0 16652 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1688980957
transform -1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1688980957
transform -1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1688980957
transform -1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1688980957
transform -1 0 16652 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1688980957
transform -1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1688980957
transform -1 0 16652 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1688980957
transform -1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1688980957
transform -1 0 16652 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1688980957
transform -1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1688980957
transform -1 0 16652 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1688980957
transform -1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1688980957
transform -1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1688980957
transform -1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1688980957
transform -1 0 16652 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1688980957
transform -1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1688980957
transform -1 0 16652 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1688980957
transform -1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1688980957
transform -1 0 16652 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1688980957
transform -1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1688980957
transform -1 0 16652 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1688980957
transform -1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_61
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_63
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_64
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_66
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_67
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_76
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_77
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_79
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_80
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_81
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_82
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_83
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_84
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_85
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_86
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_87
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_88
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_89
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_90
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_91
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_92
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_93
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_94
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_95
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_96
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_97
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_98
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_99
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_100
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_101
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_102
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_103
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_104
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_105
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_106
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_107
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_108
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_109
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_110
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_111
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_112
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_113
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_114
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_115
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_116
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_117
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_118
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_119
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_120
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_121
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_122
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_123
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_124
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_125
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_126
timestamp 1688980957
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_127
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_128
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_129
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_130
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  wb_lfsr_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
<< labels >>
flabel metal4 s 4830 2128 5150 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8717 2128 9037 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12604 2128 12924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16491 2128 16811 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2887 2128 3207 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6774 2128 7094 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10661 2128 10981 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 14548 2128 14868 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 17001 1368 17801 1488 0 FreeSans 480 0 0 0 i_clk
port 2 nsew signal input
flabel metal3 s 17001 5448 17801 5568 0 FreeSans 480 0 0 0 i_reset
port 3 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 i_wb_addr[0]
port 4 nsew signal input
flabel metal3 s 17001 13608 17801 13728 0 FreeSans 480 0 0 0 i_wb_addr[1]
port 5 nsew signal input
flabel metal3 s 17001 17688 17801 17808 0 FreeSans 480 0 0 0 i_wb_addr[2]
port 6 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 i_wb_cyc
port 7 nsew signal input
flabel metal2 s 11610 19145 11666 19945 0 FreeSans 224 90 0 0 i_wb_data[0]
port 8 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 i_wb_data[1]
port 9 nsew signal input
flabel metal2 s 3882 19145 3938 19945 0 FreeSans 224 90 0 0 i_wb_data[2]
port 10 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 i_wb_data[3]
port 11 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 i_wb_data[4]
port 12 nsew signal input
flabel metal2 s 7746 19145 7802 19945 0 FreeSans 224 90 0 0 i_wb_data[5]
port 13 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 i_wb_data[6]
port 14 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 i_wb_data[7]
port 15 nsew signal input
flabel metal2 s 15474 19145 15530 19945 0 FreeSans 224 90 0 0 i_wb_stb
port 16 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 i_wb_we
port 17 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 o_wb_ack
port 18 nsew signal tristate
flabel metal2 s 18 19145 74 19945 0 FreeSans 224 90 0 0 o_wb_data
port 19 nsew signal tristate
flabel metal3 s 17001 9528 17801 9648 0 FreeSans 480 0 0 0 o_wb_stall
port 20 nsew signal tristate
rlabel via1 8957 17408 8957 17408 0 VGND
rlabel metal1 8878 16864 8878 16864 0 VPWR
rlabel metal1 1748 12274 1748 12274 0 FLSR_instance.flip_flop_instance\[0\].in
rlabel metal2 3174 13158 3174 13158 0 FLSR_instance.flip_flop_instance\[0\].out
rlabel metal2 2346 12546 2346 12546 0 FLSR_instance.flip_flop_instance\[0\].reset
rlabel metal1 13156 15062 13156 15062 0 FLSR_instance.flip_flop_instance\[10\].in
rlabel metal2 14490 14586 14490 14586 0 FLSR_instance.flip_flop_instance\[10\].out
rlabel metal2 14398 13566 14398 13566 0 FLSR_instance.flip_flop_instance\[11\].in
rlabel metal1 14582 12954 14582 12954 0 FLSR_instance.flip_flop_instance\[11\].out
rlabel metal1 14076 11798 14076 11798 0 FLSR_instance.flip_flop_instance\[12\].in
rlabel metal1 15134 11118 15134 11118 0 FLSR_instance.flip_flop_instance\[12\].out
rlabel metal1 14950 10098 14950 10098 0 FLSR_instance.flip_flop_instance\[13\].in
rlabel metal2 14582 9792 14582 9792 0 FLSR_instance.flip_flop_instance\[13\].out
rlabel metal1 14720 9010 14720 9010 0 FLSR_instance.flip_flop_instance\[14\].in
rlabel metal1 13662 8874 13662 8874 0 FLSR_instance.flip_flop_instance\[14\].out
rlabel metal1 12512 7922 12512 7922 0 FLSR_instance.flip_flop_instance\[15\].in
rlabel metal1 14214 7786 14214 7786 0 FLSR_instance.flip_flop_instance\[15\].out
rlabel metal1 14204 6970 14204 6970 0 FLSR_instance.flip_flop_instance\[16\].in
rlabel metal1 15272 6426 15272 6426 0 FLSR_instance.flip_flop_instance\[16\].out
rlabel metal1 14444 5270 14444 5270 0 FLSR_instance.flip_flop_instance\[17\].in
rlabel metal1 15226 4590 15226 4590 0 FLSR_instance.flip_flop_instance\[17\].out
rlabel metal2 14030 4250 14030 4250 0 FLSR_instance.flip_flop_instance\[18\].in
rlabel metal1 14306 4250 14306 4250 0 FLSR_instance.flip_flop_instance\[18\].out
rlabel metal1 12236 3570 12236 3570 0 FLSR_instance.flip_flop_instance\[19\].in
rlabel metal1 13041 3366 13041 3366 0 FLSR_instance.flip_flop_instance\[19\].out
rlabel metal1 2622 12920 2622 12920 0 FLSR_instance.flip_flop_instance\[1\].in
rlabel metal2 4738 13634 4738 13634 0 FLSR_instance.flip_flop_instance\[1\].out
rlabel metal1 10028 4182 10028 4182 0 FLSR_instance.flip_flop_instance\[20\].in
rlabel metal1 11776 4046 11776 4046 0 FLSR_instance.flip_flop_instance\[20\].out
rlabel metal1 10488 5338 10488 5338 0 FLSR_instance.flip_flop_instance\[21\].in
rlabel metal1 9936 5610 9936 5610 0 FLSR_instance.flip_flop_instance\[21\].out
rlabel metal1 8004 5746 8004 5746 0 FLSR_instance.flip_flop_instance\[22\].in
rlabel metal1 9062 5814 9062 5814 0 FLSR_instance.flip_flop_instance\[22\].out
rlabel metal1 6440 5882 6440 5882 0 FLSR_instance.flip_flop_instance\[23\].in
rlabel metal1 7728 6426 7728 6426 0 FLSR_instance.flip_flop_instance\[23\].out
rlabel metal1 3128 5270 3128 5270 0 FLSR_instance.flip_flop_instance\[24\].in
rlabel metal2 4186 4250 4186 4250 0 FLSR_instance.flip_flop_instance\[24\].out
rlabel metal1 3772 4182 3772 4182 0 FLSR_instance.flip_flop_instance\[25\].in
rlabel metal2 5198 4420 5198 4420 0 FLSR_instance.flip_flop_instance\[25\].out
rlabel metal1 5704 4658 5704 4658 0 FLSR_instance.flip_flop_instance\[26\].in
rlabel metal1 7360 3502 7360 3502 0 FLSR_instance.flip_flop_instance\[26\].out
rlabel metal1 6946 4046 6946 4046 0 FLSR_instance.flip_flop_instance\[27\].in
rlabel metal1 7084 4250 7084 4250 0 FLSR_instance.flip_flop_instance\[27\].out
rlabel metal1 4692 5882 4692 5882 0 FLSR_instance.flip_flop_instance\[28\].in
rlabel metal1 5888 6154 5888 6154 0 FLSR_instance.flip_flop_instance\[28\].out
rlabel metal1 3680 6970 3680 6970 0 FLSR_instance.flip_flop_instance\[29\].in
rlabel metal1 4554 7514 4554 7514 0 FLSR_instance.flip_flop_instance\[29\].out
rlabel metal1 5842 14450 5842 14450 0 FLSR_instance.flip_flop_instance\[2\].in
rlabel metal1 7590 14586 7590 14586 0 FLSR_instance.flip_flop_instance\[2\].out
rlabel metal1 2898 8058 2898 8058 0 FLSR_instance.flip_flop_instance\[30\].in
rlabel metal1 4140 8602 4140 8602 0 FLSR_instance.flip_flop_instance\[30\].out
rlabel metal1 3772 9962 3772 9962 0 FLSR_instance.flip_flop_instance\[31\].in
rlabel metal2 5566 11254 5566 11254 0 FLSR_instance.flip_flop_instance\[31\].out
rlabel metal1 7406 16218 7406 16218 0 FLSR_instance.flip_flop_instance\[3\].in
rlabel metal1 9062 16762 9062 16762 0 FLSR_instance.flip_flop_instance\[3\].out
rlabel metal2 6486 16422 6486 16422 0 FLSR_instance.flip_flop_instance\[4\].in
rlabel metal1 7038 16762 7038 16762 0 FLSR_instance.flip_flop_instance\[4\].out
rlabel metal1 5014 15674 5014 15674 0 FLSR_instance.flip_flop_instance\[5\].in
rlabel metal1 6026 12954 6026 12954 0 FLSR_instance.flip_flop_instance\[5\].out
rlabel metal1 6210 12410 6210 12410 0 FLSR_instance.flip_flop_instance\[6\].in
rlabel metal1 6256 12070 6256 12070 0 FLSR_instance.flip_flop_instance\[6\].out
rlabel metal1 8602 13226 8602 13226 0 FLSR_instance.flip_flop_instance\[7\].in
rlabel metal1 10534 13498 10534 13498 0 FLSR_instance.flip_flop_instance\[7\].out
rlabel metal1 9844 14586 9844 14586 0 FLSR_instance.flip_flop_instance\[8\].in
rlabel metal1 11638 15130 11638 15130 0 FLSR_instance.flip_flop_instance\[8\].out
rlabel metal1 11500 16150 11500 16150 0 FLSR_instance.flip_flop_instance\[9\].in
rlabel metal1 13524 16218 13524 16218 0 FLSR_instance.flip_flop_instance\[9\].out
rlabel metal1 5014 13804 5014 13804 0 FLSR_instance.load_seed
rlabel metal1 2898 16082 2898 16082 0 FLSR_instance.muxes\[0\].input_a
rlabel metal2 13202 15300 13202 15300 0 FLSR_instance.muxes\[10\].input_a
rlabel metal2 14306 13464 14306 13464 0 FLSR_instance.muxes\[11\].input_a
rlabel metal1 13524 12410 13524 12410 0 FLSR_instance.muxes\[12\].input_a
rlabel metal1 13662 11220 13662 11220 0 FLSR_instance.muxes\[13\].input_a
rlabel metal1 14306 9622 14306 9622 0 FLSR_instance.muxes\[14\].input_a
rlabel metal1 12880 9418 12880 9418 0 FLSR_instance.muxes\[15\].input_a
rlabel metal1 13386 7480 13386 7480 0 FLSR_instance.muxes\[16\].input_a
rlabel metal1 14260 6154 14260 6154 0 FLSR_instance.muxes\[17\].input_a
rlabel metal1 14122 4658 14122 4658 0 FLSR_instance.muxes\[18\].input_a
rlabel metal1 12742 2346 12742 2346 0 FLSR_instance.muxes\[19\].input_a
rlabel metal1 3266 13158 3266 13158 0 FLSR_instance.muxes\[1\].input_a
rlabel metal1 10350 2346 10350 2346 0 FLSR_instance.muxes\[20\].input_a
rlabel metal1 11408 7174 11408 7174 0 FLSR_instance.muxes\[21\].input_a
rlabel metal1 9844 5338 9844 5338 0 FLSR_instance.muxes\[22\].input_a
rlabel metal2 9890 6970 9890 6970 0 FLSR_instance.muxes\[23\].input_a
rlabel metal2 7406 7616 7406 7616 0 FLSR_instance.muxes\[24\].input_a
rlabel metal1 3542 2346 3542 2346 0 FLSR_instance.muxes\[25\].input_a
rlabel metal1 3128 4726 3128 4726 0 FLSR_instance.muxes\[26\].input_a
rlabel metal1 7682 3162 7682 3162 0 FLSR_instance.muxes\[27\].input_a
rlabel metal1 5520 2346 5520 2346 0 FLSR_instance.muxes\[28\].input_a
rlabel metal1 5980 7854 5980 7854 0 FLSR_instance.muxes\[29\].input_a
rlabel metal1 5014 14042 5014 14042 0 FLSR_instance.muxes\[2\].input_a
rlabel metal1 2484 6766 2484 6766 0 FLSR_instance.muxes\[30\].input_a
rlabel metal1 2507 8942 2507 8942 0 FLSR_instance.muxes\[31\].input_a
rlabel metal1 8740 14042 8740 14042 0 FLSR_instance.muxes\[3\].input_a
rlabel metal1 9384 16218 9384 16218 0 FLSR_instance.muxes\[4\].input_a
rlabel metal1 5474 17306 5474 17306 0 FLSR_instance.muxes\[5\].input_a
rlabel metal2 5934 12585 5934 12585 0 FLSR_instance.muxes\[6\].input_a
rlabel metal2 7958 11322 7958 11322 0 FLSR_instance.muxes\[7\].input_a
rlabel metal2 11086 13396 11086 13396 0 FLSR_instance.muxes\[8\].input_a
rlabel metal1 12098 12410 12098 12410 0 FLSR_instance.muxes\[9\].input_a
rlabel metal2 4554 9826 4554 9826 0 _000_
rlabel metal2 4002 8636 4002 8636 0 _001_
rlabel metal1 4883 7446 4883 7446 0 _002_
rlabel metal1 5336 5882 5336 5882 0 _003_
rlabel metal2 7774 4318 7774 4318 0 _004_
rlabel metal1 7275 4522 7275 4522 0 _005_
rlabel metal2 4462 4318 4462 4318 0 _006_
rlabel metal2 4002 5406 4002 5406 0 _007_
rlabel metal1 6992 5882 6992 5882 0 _008_
rlabel metal1 8142 5338 8142 5338 0 _009_
rlabel metal1 12289 5610 12289 5610 0 _010_
rlabel metal1 11638 4148 11638 4148 0 _011_
rlabel metal1 13623 3434 13623 3434 0 _012_
rlabel metal1 15686 4148 15686 4148 0 _013_
rlabel metal1 15923 5270 15923 5270 0 _014_
rlabel metal1 15272 7174 15272 7174 0 _015_
rlabel metal2 13754 7650 13754 7650 0 _016_
rlabel metal1 15831 8874 15831 8874 0 _017_
rlabel metal2 15410 9826 15410 9826 0 _018_
rlabel metal1 14996 10778 14996 10778 0 _019_
rlabel metal1 14950 13974 14950 13974 0 _020_
rlabel metal2 14214 15198 14214 15198 0 _021_
rlabel metal2 12282 15912 12282 15912 0 _022_
rlabel metal1 10626 14586 10626 14586 0 _023_
rlabel metal2 9522 13090 9522 13090 0 _024_
rlabel metal1 7038 12410 7038 12410 0 _025_
rlabel metal2 6302 15912 6302 15912 0 _026_
rlabel metal1 6900 16218 6900 16218 0 _027_
rlabel metal2 8418 16388 8418 16388 0 _028_
rlabel metal1 7367 14314 7367 14314 0 _029_
rlabel metal1 4094 12410 4094 12410 0 _030_
rlabel metal1 2806 12648 2806 12648 0 _031_
rlabel metal1 6706 7854 6706 7854 0 _032_
rlabel metal1 2806 3128 2806 3128 0 _033_
rlabel via1 1697 4590 1697 4590 0 _034_
rlabel metal1 7084 2618 7084 2618 0 _035_
rlabel via1 4728 3094 4728 3094 0 _036_
rlabel metal1 5147 8534 5147 8534 0 _037_
rlabel metal2 1702 7174 1702 7174 0 _038_
rlabel metal1 1656 9146 1656 9146 0 _039_
rlabel metal1 12174 7446 12174 7446 0 _040_
rlabel metal1 12519 6358 12519 6358 0 _041_
rlabel metal1 12473 5270 12473 5270 0 _042_
rlabel metal1 12328 2618 12328 2618 0 _043_
rlabel metal1 10299 3026 10299 3026 0 _044_
rlabel metal2 11086 7174 11086 7174 0 _045_
rlabel metal2 9798 4998 9798 4998 0 _046_
rlabel metal1 9517 7446 9517 7446 0 _047_
rlabel metal2 6946 9826 6946 9826 0 _048_
rlabel metal2 2162 16354 2162 16354 0 _049_
rlabel via1 2249 11118 2249 11118 0 _050_
rlabel metal1 3526 14314 3526 14314 0 _051_
rlabel metal1 7815 13974 7815 13974 0 _052_
rlabel metal2 9798 16354 9798 16354 0 _053_
rlabel metal2 3910 16966 3910 16966 0 _054_
rlabel metal1 4876 10778 4876 10778 0 _055_
rlabel metal1 6762 10778 6762 10778 0 _056_
rlabel metal2 11362 13090 11362 13090 0 _057_
rlabel metal2 12098 12002 12098 12002 0 _058_
rlabel metal2 12374 14178 12374 14178 0 _059_
rlabel metal1 12972 13498 12972 13498 0 _060_
rlabel via1 12553 12206 12553 12206 0 _061_
rlabel metal1 12374 11152 12374 11152 0 _062_
rlabel metal1 12634 9962 12634 9962 0 _063_
rlabel metal1 11582 9554 11582 9554 0 _064_
rlabel via1 1697 10710 1697 10710 0 _065_
rlabel metal2 1702 14790 1702 14790 0 _066_
rlabel metal1 9292 11866 9292 11866 0 _067_
rlabel metal1 5842 4012 5842 4012 0 _068_
rlabel metal1 3588 9690 3588 9690 0 _069_
rlabel metal1 3496 7854 3496 7854 0 _070_
rlabel metal1 4692 6766 4692 6766 0 _071_
rlabel metal2 5290 4301 5290 4301 0 _072_
rlabel metal1 6854 3706 6854 3706 0 _073_
rlabel metal2 4738 4998 4738 4998 0 _074_
rlabel metal1 3910 3706 3910 3706 0 _075_
rlabel metal1 3450 6358 3450 6358 0 _076_
rlabel metal1 6394 5644 6394 5644 0 _077_
rlabel metal1 14904 9486 14904 9486 0 _078_
rlabel metal1 9016 5882 9016 5882 0 _079_
rlabel metal1 10718 5236 10718 5236 0 _080_
rlabel metal2 10350 4148 10350 4148 0 _081_
rlabel metal1 12650 4114 12650 4114 0 _082_
rlabel metal1 14030 4590 14030 4590 0 _083_
rlabel metal1 14444 5678 14444 5678 0 _084_
rlabel metal1 14168 7378 14168 7378 0 _085_
rlabel metal1 12742 8466 12742 8466 0 _086_
rlabel metal1 14720 9554 14720 9554 0 _087_
rlabel metal1 15272 10642 15272 10642 0 _088_
rlabel metal1 14214 14450 14214 14450 0 _089_
rlabel metal1 13386 12614 13386 12614 0 _090_
rlabel metal1 14858 13872 14858 13872 0 _091_
rlabel metal1 13202 15470 13202 15470 0 _092_
rlabel metal1 11454 14858 11454 14858 0 _093_
rlabel metal2 9982 14212 9982 14212 0 _094_
rlabel metal1 7728 13294 7728 13294 0 _095_
rlabel metal1 5612 12614 5612 12614 0 _096_
rlabel metal1 5382 15470 5382 15470 0 _097_
rlabel metal1 6670 16116 6670 16116 0 _098_
rlabel metal1 7544 15130 7544 15130 0 _099_
rlabel metal1 4554 14042 4554 14042 0 _100_
rlabel metal2 2714 12988 2714 12988 0 _101_
rlabel metal1 5290 12410 5290 12410 0 _102_
rlabel metal1 5198 13498 5198 13498 0 _103_
rlabel metal1 2530 14246 2530 14246 0 _104_
rlabel metal1 2162 13906 2162 13906 0 _105_
rlabel metal1 2392 8466 2392 8466 0 _106_
rlabel metal1 7912 7514 7912 7514 0 _107_
rlabel metal1 8280 10642 8280 10642 0 _108_
rlabel metal1 8372 8806 8372 8806 0 _109_
rlabel metal1 9246 9010 9246 9010 0 _110_
rlabel metal1 3772 2482 3772 2482 0 _111_
rlabel metal1 7084 7514 7084 7514 0 _112_
rlabel metal1 3818 2414 3818 2414 0 _113_
rlabel metal1 2852 2618 2852 2618 0 _114_
rlabel metal2 3082 5440 3082 5440 0 _115_
rlabel metal1 1840 5202 1840 5202 0 _116_
rlabel metal1 8786 3094 8786 3094 0 _117_
rlabel metal1 7222 2448 7222 2448 0 _118_
rlabel metal2 5382 2587 5382 2587 0 _119_
rlabel metal1 4830 2618 4830 2618 0 _120_
rlabel metal2 5842 8364 5842 8364 0 _121_
rlabel metal2 5382 8500 5382 8500 0 _122_
rlabel metal1 2806 6630 2806 6630 0 _123_
rlabel metal1 1932 6630 1932 6630 0 _124_
rlabel metal1 2392 8602 2392 8602 0 _125_
rlabel metal1 1840 8942 1840 8942 0 _126_
rlabel metal1 10718 8500 10718 8500 0 _127_
rlabel metal1 10764 10642 10764 10642 0 _128_
rlabel metal1 12052 2414 12052 2414 0 _129_
rlabel metal1 11178 9112 11178 9112 0 _130_
rlabel metal1 10902 7888 10902 7888 0 _131_
rlabel metal1 10166 2312 10166 2312 0 _132_
rlabel metal1 8234 9146 8234 9146 0 _133_
rlabel metal1 8188 9622 8188 9622 0 _134_
rlabel metal1 8510 10574 8510 10574 0 _135_
rlabel metal1 7314 9554 7314 9554 0 _136_
rlabel metal1 3588 14382 3588 14382 0 _137_
rlabel metal1 3450 16150 3450 16150 0 _138_
rlabel metal1 3266 15980 3266 15980 0 _139_
rlabel metal1 2484 16082 2484 16082 0 _140_
rlabel metal1 3358 10676 3358 10676 0 _141_
rlabel metal1 2852 10778 2852 10778 0 _142_
rlabel metal1 3772 14042 3772 14042 0 _143_
rlabel metal1 3312 14042 3312 14042 0 _144_
rlabel metal1 9384 14042 9384 14042 0 _145_
rlabel metal1 8510 14382 8510 14382 0 _146_
rlabel metal2 9430 15844 9430 15844 0 _147_
rlabel metal1 9982 16014 9982 16014 0 _148_
rlabel metal2 5198 16014 5198 16014 0 _149_
rlabel metal1 4186 16558 4186 16558 0 _150_
rlabel metal2 5842 10914 5842 10914 0 _151_
rlabel metal1 5198 10676 5198 10676 0 _152_
rlabel metal2 7498 10880 7498 10880 0 _153_
rlabel metal1 7038 10710 7038 10710 0 _154_
rlabel metal1 11362 9146 11362 9146 0 _155_
rlabel metal1 12604 13294 12604 13294 0 _156_
rlabel metal1 11408 10642 11408 10642 0 _157_
rlabel metal1 12558 13192 12558 13192 0 _158_
rlabel metal1 1886 11662 1886 11662 0 _159_
rlabel metal1 2622 14518 2622 14518 0 _160_
rlabel metal1 1932 14382 1932 14382 0 _161_
rlabel metal2 9982 10642 9982 10642 0 _162_
rlabel metal1 9292 11322 9292 11322 0 _163_
rlabel metal1 4462 9588 4462 9588 0 _164_
rlabel metal1 14858 10676 14858 10676 0 _165_
rlabel metal1 14398 13974 14398 13974 0 _166_
rlabel metal1 16376 2414 16376 2414 0 i_clk
rlabel metal1 16652 5678 16652 5678 0 i_reset
rlabel metal2 11638 823 11638 823 0 i_wb_addr[0]
rlabel metal1 16330 13906 16330 13906 0 i_wb_addr[1]
rlabel metal2 15962 17493 15962 17493 0 i_wb_addr[2]
rlabel metal3 820 16388 820 16388 0 i_wb_cyc
rlabel metal1 11730 17238 11730 17238 0 i_wb_data[0]
rlabel metal2 46 1588 46 1588 0 i_wb_data[1]
rlabel metal1 3542 17238 3542 17238 0 i_wb_data[2]
rlabel metal2 15502 959 15502 959 0 i_wb_data[3]
rlabel metal2 3910 959 3910 959 0 i_wb_data[4]
rlabel metal1 7866 17238 7866 17238 0 i_wb_data[5]
rlabel metal3 820 4148 820 4148 0 i_wb_data[6]
rlabel metal3 1050 8228 1050 8228 0 i_wb_data[7]
rlabel metal1 15548 17170 15548 17170 0 i_wb_stb
rlabel metal2 7774 1588 7774 1588 0 i_wb_we
rlabel metal1 15134 3434 15134 3434 0 net1
rlabel metal1 11822 2482 11822 2482 0 net10
rlabel metal1 5014 2278 5014 2278 0 net11
rlabel metal3 7682 12716 7682 12716 0 net12
rlabel metal2 2714 4760 2714 4760 0 net13
rlabel metal1 2070 8364 2070 8364 0 net14
rlabel metal2 15778 11696 15778 11696 0 net15
rlabel metal1 8234 2618 8234 2618 0 net16
rlabel metal1 1518 12784 1518 12784 0 net17
rlabel metal2 2346 14756 2346 14756 0 net18
rlabel metal1 6578 2618 6578 2618 0 net19
rlabel metal2 16146 8466 16146 8466 0 net2
rlabel metal1 1472 7378 1472 7378 0 net20
rlabel metal1 13754 4148 13754 4148 0 net21
rlabel metal2 13938 7888 13938 7888 0 net22
rlabel metal1 1702 16694 1702 16694 0 net23
rlabel metal1 3450 14450 3450 14450 0 net24
rlabel metal1 12512 10098 12512 10098 0 net25
rlabel metal1 13984 13362 13984 13362 0 net26
rlabel metal1 6532 2414 6532 2414 0 net27
rlabel via2 16330 9571 16330 9571 0 net28
rlabel metal1 12558 2618 12558 2618 0 net3
rlabel metal1 12466 14280 12466 14280 0 net4
rlabel metal1 16054 17000 16054 17000 0 net5
rlabel metal1 2162 16422 2162 16422 0 net6
rlabel metal2 11914 16286 11914 16286 0 net7
rlabel metal1 2760 2550 2760 2550 0 net8
rlabel metal1 11684 13906 11684 13906 0 net9
rlabel metal3 1142 12308 1142 12308 0 o_wb_ack
rlabel metal1 828 17306 828 17306 0 o_wb_data
<< properties >>
string FIXED_BBOX 0 0 17801 19945
<< end >>
