magic
tech sky130A
magscale 1 2
timestamp 1692995762
<< obsli1 >>
rect 1104 2159 16652 17425
<< obsm1 >>
rect 14 2128 17006 17456
<< metal2 >>
rect 18 19145 74 19945
rect 3882 19145 3938 19945
rect 7746 19145 7802 19945
rect 11610 19145 11666 19945
rect 15474 19145 15530 19945
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 15474 0 15530 800
<< obsm2 >>
rect 130 19089 3826 19258
rect 3994 19089 7690 19258
rect 7858 19089 11554 19258
rect 11722 19089 15418 19258
rect 15586 19089 17002 19258
rect 20 856 17002 19089
rect 130 734 3826 856
rect 3994 734 7690 856
rect 7858 734 11554 856
rect 11722 734 15418 856
rect 15586 734 17002 856
<< metal3 >>
rect 17001 17688 17801 17808
rect 0 16328 800 16448
rect 17001 13608 17801 13728
rect 0 12248 800 12368
rect 17001 9528 17801 9648
rect 0 8168 800 8288
rect 17001 5448 17801 5568
rect 0 4088 800 4208
rect 17001 1368 17801 1488
<< obsm3 >>
rect 800 17608 16921 17781
rect 800 16528 17001 17608
rect 880 16248 17001 16528
rect 800 13808 17001 16248
rect 800 13528 16921 13808
rect 800 12448 17001 13528
rect 880 12168 17001 12448
rect 800 9728 17001 12168
rect 800 9448 16921 9728
rect 800 8368 17001 9448
rect 880 8088 17001 8368
rect 800 5648 17001 8088
rect 800 5368 16921 5648
rect 800 4288 17001 5368
rect 880 4008 17001 4288
rect 800 1568 17001 4008
rect 800 1395 16921 1568
<< metal4 >>
rect 2887 2128 3207 17456
rect 4830 2128 5150 17456
rect 6774 2128 7094 17456
rect 8717 2128 9037 17456
rect 10661 2128 10981 17456
rect 12604 2128 12924 17456
rect 14548 2128 14868 17456
rect 16491 2128 16811 17456
<< labels >>
rlabel metal4 s 4830 2128 5150 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8717 2128 9037 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 16491 2128 16811 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2887 2128 3207 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6774 2128 7094 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 10661 2128 10981 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 14548 2128 14868 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 17001 1368 17801 1488 6 i_clk
port 3 nsew signal input
rlabel metal3 s 17001 5448 17801 5568 6 i_reset
port 4 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 i_wb_addr[0]
port 5 nsew signal input
rlabel metal3 s 17001 13608 17801 13728 6 i_wb_addr[1]
port 6 nsew signal input
rlabel metal3 s 17001 17688 17801 17808 6 i_wb_addr[2]
port 7 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 i_wb_cyc
port 8 nsew signal input
rlabel metal2 s 11610 19145 11666 19945 6 i_wb_data[0]
port 9 nsew signal input
rlabel metal2 s 18 0 74 800 6 i_wb_data[1]
port 10 nsew signal input
rlabel metal2 s 3882 19145 3938 19945 6 i_wb_data[2]
port 11 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 i_wb_data[3]
port 12 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 i_wb_data[4]
port 13 nsew signal input
rlabel metal2 s 7746 19145 7802 19945 6 i_wb_data[5]
port 14 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 i_wb_data[6]
port 15 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 i_wb_data[7]
port 16 nsew signal input
rlabel metal2 s 15474 19145 15530 19945 6 i_wb_stb
port 17 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 i_wb_we
port 18 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 o_wb_ack
port 19 nsew signal output
rlabel metal2 s 18 19145 74 19945 6 o_wb_data
port 20 nsew signal output
rlabel metal3 s 17001 9528 17801 9648 6 o_wb_stall
port 21 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 17801 19945
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 915288
string GDS_FILE /openlane/designs/wb_lfsr/runs/RUN_2023.08.25_20.34.39/results/signoff/wb_lfsr.magic.gds
string GDS_START 229646
<< end >>

