* NGSPICE file created from wb_lfsr.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt wb_lfsr VGND VPWR i_clk i_reset i_wb_addr[0] i_wb_addr[1] i_wb_addr[2] i_wb_cyc
+ i_wb_data[0] i_wb_data[1] i_wb_data[2] i_wb_data[3] i_wb_data[4] i_wb_data[5] i_wb_data[6]
+ i_wb_data[7] i_wb_stb i_wb_we o_wb_ack o_wb_data o_wb_stall
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_363_ _166_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
X_294_ FLSR_instance.muxes\[2\].input_a _143_ _139_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__mux2_1
X_432_ net23 FLSR_instance.flip_flop_instance\[1\].in _030_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[1\].out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_415_ net21 FLSR_instance.flip_flop_instance\[18\].in _013_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[18\].out
+ sky130_fd_sc_hd__dfrtp_1
X_346_ _165_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__inv_2
X_277_ FLSR_instance.muxes\[21\].input_a _129_ _132_ net12 VGND VGND VPWR VPWR _045_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_200_ _085_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[16\].in sky130_fd_sc_hd__clkbuf_1
X_329_ FLSR_instance.flip_flop_instance\[0\].reset _162_ _135_ VGND VGND VPWR VPWR
+ _163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_362_ _166_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_431_ net24 FLSR_instance.flip_flop_instance\[2\].in _029_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[2\].out
+ sky130_fd_sc_hd__dfrtp_1
X_293_ net9 _137_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_21_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _165_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__inv_2
X_414_ net21 FLSR_instance.flip_flop_instance\[19\].in _012_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[19\].out
+ sky130_fd_sc_hd__dfrtp_1
X_276_ FLSR_instance.muxes\[20\].input_a _129_ _132_ net11 VGND VGND VPWR VPWR _044_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_328_ net7 net4 net3 VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__or3_1
X_259_ _122_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_24_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_430_ net24 FLSR_instance.flip_flop_instance\[3\].in _028_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[3\].out
+ sky130_fd_sc_hd__dfrtp_1
X_361_ _166_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__inv_2
X_292_ _142_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_275_ FLSR_instance.muxes\[19\].input_a _129_ _132_ net10 VGND VGND VPWR VPWR _043_
+ sky130_fd_sc_hd__a22o_1
X_413_ net21 FLSR_instance.flip_flop_instance\[20\].in _011_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[20\].out
+ sky130_fd_sc_hd__dfrtp_1
X_344_ _165_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_327_ _161_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__clkbuf_1
X_189_ FLSR_instance.flip_flop_instance\[20\].out FLSR_instance.muxes\[21\].input_a
+ _078_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__mux2_1
X_258_ FLSR_instance.muxes\[29\].input_a _121_ _111_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _166_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__inv_2
X_291_ FLSR_instance.muxes\[1\].input_a _141_ _139_ VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_274_ FLSR_instance.muxes\[18\].input_a _129_ _132_ net9 VGND VGND VPWR VPWR _042_
+ sky130_fd_sc_hd__a22o_1
X_412_ net21 FLSR_instance.flip_flop_instance\[21\].in _010_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[21\].out
+ sky130_fd_sc_hd__dfrtp_1
X_343_ _165_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_326_ net18 _104_ _160_ VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__mux2_1
X_188_ _079_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[22\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_257_ net12 _106_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_309_ FLSR_instance.muxes\[7\].input_a _153_ _139_ VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_290_ net8 _137_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_342_ FLSR_instance.flip_flop_instance\[0\].reset VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__buf_4
X_411_ net19 FLSR_instance.flip_flop_instance\[22\].in _009_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[22\].out
+ sky130_fd_sc_hd__dfrtp_1
X_273_ FLSR_instance.muxes\[17\].input_a _129_ _132_ net8 VGND VGND VPWR VPWR _041_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_325_ net16 net6 net15 VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__and3b_1
X_256_ _120_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_187_ FLSR_instance.flip_flop_instance\[21\].out FLSR_instance.muxes\[22\].input_a
+ _078_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_239_ net15 net16 net6 VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__and3_1
X_308_ net14 _137_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_341_ _164_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
X_410_ net20 FLSR_instance.flip_flop_instance\[23\].in _008_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[23\].out
+ sky130_fd_sc_hd__dfrtp_1
X_272_ FLSR_instance.muxes\[16\].input_a _129_ _132_ net7 VGND VGND VPWR VPWR _040_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_324_ _159_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__clkbuf_1
X_186_ FLSR_instance.load_seed VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_13_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_255_ FLSR_instance.muxes\[28\].input_a _119_ _111_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_307_ _152_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__clkbuf_1
X_169_ _069_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[31\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_238_ net7 _106_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_340_ _164_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__inv_2
X_271_ _131_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__buf_2
X_323_ net2 net15 VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_13_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_254_ net11 _106_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__and2_1
X_185_ _077_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[23\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_306_ FLSR_instance.muxes\[6\].input_a _151_ _139_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__mux2_1
X_168_ FLSR_instance.flip_flop_instance\[30\].out FLSR_instance.muxes\[31\].input_a
+ _068_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__mux2_1
X_237_ net5 net4 net3 VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__and3b_2
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_270_ _127_ _130_ _128_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__and3_1
X_399_ net23 _065_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_1
X_322_ FLSR_instance.muxes\[15\].input_a _156_ _158_ net14 VGND VGND VPWR VPWR _064_
+ sky130_fd_sc_hd__a22o_1
X_253_ _118_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__clkbuf_1
X_184_ FLSR_instance.flip_flop_instance\[22\].out FLSR_instance.muxes\[23\].input_a
+ _068_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_236_ _105_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[0\].in sky130_fd_sc_hd__clkbuf_1
X_305_ net13 _137_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__and2_1
X_167_ FLSR_instance.load_seed VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_219_ _095_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[7\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_398_ net22 _064_ VGND VGND VPWR VPWR FLSR_instance.muxes\[15\].input_a sky130_fd_sc_hd__dfxtp_1
X_321_ FLSR_instance.muxes\[14\].input_a _156_ _158_ net13 VGND VGND VPWR VPWR _063_
+ sky130_fd_sc_hd__a22o_1
X_252_ FLSR_instance.muxes\[27\].input_a _117_ _111_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__mux2_1
X_183_ _076_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[24\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_304_ _150_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__clkbuf_1
X_235_ _104_ FLSR_instance.muxes\[0\].input_a FLSR_instance.load_seed VGND VGND VPWR
+ VPWR _105_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_7_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_218_ FLSR_instance.flip_flop_instance\[6\].out FLSR_instance.muxes\[7\].input_a
+ _089_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput17 net17 VGND VGND VPWR VPWR o_wb_ack sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_397_ net25 _063_ VGND VGND VPWR VPWR FLSR_instance.muxes\[14\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_320_ FLSR_instance.muxes\[13\].input_a _156_ _158_ net12 VGND VGND VPWR VPWR _062_
+ sky130_fd_sc_hd__a22o_1
X_251_ net10 _106_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__and2_1
X_182_ FLSR_instance.flip_flop_instance\[23\].out FLSR_instance.muxes\[24\].input_a
+ _068_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_303_ FLSR_instance.muxes\[5\].input_a _149_ _139_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_23_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_234_ _102_ _103_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_10_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_217_ _094_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[8\].in sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput18 net18 VGND VGND VPWR VPWR o_wb_data sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_26_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_396_ net25 _062_ VGND VGND VPWR VPWR FLSR_instance.muxes\[13\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_181_ _075_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[25\].in sky130_fd_sc_hd__clkbuf_1
X_250_ _116_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__clkbuf_1
Xfanout20 net27 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_379_ net22 _045_ VGND VGND VPWR VPWR FLSR_instance.muxes\[21\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_302_ net12 _137_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__and2_1
X_233_ FLSR_instance.flip_flop_instance\[5\].out FLSR_instance.flip_flop_instance\[1\].out
+ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_216_ FLSR_instance.flip_flop_instance\[7\].out FLSR_instance.muxes\[8\].input_a
+ _089_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_395_ net25 _061_ VGND VGND VPWR VPWR FLSR_instance.muxes\[12\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout21 net27 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
X_180_ FLSR_instance.flip_flop_instance\[24\].out FLSR_instance.muxes\[25\].input_a
+ _068_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_378_ net21 _044_ VGND VGND VPWR VPWR FLSR_instance.muxes\[20\].input_a sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_301_ _148_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__clkbuf_1
X_232_ FLSR_instance.flip_flop_instance\[6\].out FLSR_instance.flip_flop_instance\[31\].out
+ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_215_ _093_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[9\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_394_ net26 _060_ VGND VGND VPWR VPWR FLSR_instance.muxes\[11\].input_a sky130_fd_sc_hd__dfxtp_1
Xfanout22 net27 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
X_377_ net21 _043_ VGND VGND VPWR VPWR FLSR_instance.muxes\[19\].input_a sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_300_ FLSR_instance.muxes\[4\].input_a _147_ _139_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_231_ _101_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[1\].in sky130_fd_sc_hd__clkbuf_1
X_429_ net24 FLSR_instance.flip_flop_instance\[4\].in _027_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[4\].out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput1 i_clk VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_214_ FLSR_instance.flip_flop_instance\[8\].out FLSR_instance.muxes\[9\].input_a
+ _089_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_393_ net25 _059_ VGND VGND VPWR VPWR FLSR_instance.muxes\[10\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout23 net27 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ net21 _042_ VGND VGND VPWR VPWR FLSR_instance.muxes\[18\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_230_ FLSR_instance.flip_flop_instance\[0\].out FLSR_instance.muxes\[1\].input_a
+ FLSR_instance.load_seed VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__mux2_1
X_428_ net24 FLSR_instance.flip_flop_instance\[5\].in _026_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[5\].out
+ sky130_fd_sc_hd__dfrtp_1
X_359_ _166_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 i_reset VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_213_ _092_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[10\].in sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_392_ net25 _058_ VGND VGND VPWR VPWR FLSR_instance.muxes\[9\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout24 net27 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_375_ net22 _041_ VGND VGND VPWR VPWR FLSR_instance.muxes\[17\].input_a sky130_fd_sc_hd__dfxtp_1
X_358_ _166_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__inv_2
X_427_ net23 FLSR_instance.flip_flop_instance\[6\].in _025_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[6\].out
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ _140_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 i_wb_addr[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_212_ FLSR_instance.flip_flop_instance\[9\].out FLSR_instance.muxes\[10\].input_a
+ _089_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_391_ net25 _057_ VGND VGND VPWR VPWR FLSR_instance.muxes\[8\].input_a sky130_fd_sc_hd__dfxtp_1
Xfanout25 net27 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_374_ net21 _040_ VGND VGND VPWR VPWR FLSR_instance.muxes\[16\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_288_ FLSR_instance.muxes\[0\].input_a _138_ _139_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__mux2_1
X_357_ _166_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__inv_2
Xinput4 i_wb_addr[1] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
X_426_ net26 FLSR_instance.flip_flop_instance\[7\].in _024_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[7\].out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_211_ _091_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[11\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_409_ net19 FLSR_instance.flip_flop_instance\[24\].in _007_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[24\].out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_390_ net23 _056_ VGND VGND VPWR VPWR FLSR_instance.muxes\[7\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout26 net27 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_18_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_373_ net20 _039_ VGND VGND VPWR VPWR FLSR_instance.muxes\[31\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 i_wb_addr[2] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_4
X_356_ _166_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_425_ net26 FLSR_instance.flip_flop_instance\[8\].in _023_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[8\].out
+ sky130_fd_sc_hd__dfrtp_1
X_287_ net5 _127_ _108_ _109_ _110_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__o2111a_4
X_210_ FLSR_instance.flip_flop_instance\[10\].out FLSR_instance.muxes\[11\].input_a
+ _089_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__mux2_1
X_408_ net19 FLSR_instance.flip_flop_instance\[25\].in _006_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[25\].out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_339_ _164_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout27 net1 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
X_372_ net20 _038_ VGND VGND VPWR VPWR FLSR_instance.muxes\[30\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_424_ net26 FLSR_instance.flip_flop_instance\[9\].in _022_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[9\].out
+ sky130_fd_sc_hd__dfrtp_1
X_286_ net7 _137_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__and2_1
X_355_ _166_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 i_wb_cyc VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ _164_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__inv_2
X_407_ net19 FLSR_instance.flip_flop_instance\[26\].in _005_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[26\].out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_269_ net5 net4 VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_25_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_371_ net20 _037_ VGND VGND VPWR VPWR FLSR_instance.muxes\[29\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_423_ net26 FLSR_instance.flip_flop_instance\[10\].in _021_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[10\].out
+ sky130_fd_sc_hd__dfrtp_1
X_354_ _166_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__inv_2
X_285_ net5 net4 net3 VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__nor3_2
XFILLER_0_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 i_wb_data[0] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_1_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_406_ net19 FLSR_instance.flip_flop_instance\[27\].in _004_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[27\].out
+ sky130_fd_sc_hd__dfrtp_1
X_337_ _164_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__inv_2
X_199_ FLSR_instance.flip_flop_instance\[15\].out FLSR_instance.muxes\[16\].input_a
+ _078_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__mux2_1
X_268_ net5 _127_ _128_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_25_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 i_wb_data[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_370_ net19 _036_ VGND VGND VPWR VPWR FLSR_instance.muxes\[28\].input_a sky130_fd_sc_hd__dfxtp_1
X_422_ net26 FLSR_instance.flip_flop_instance\[11\].in _020_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[11\].out
+ sky130_fd_sc_hd__dfrtp_1
X_353_ FLSR_instance.flip_flop_instance\[0\].reset VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_284_ _136_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 i_wb_data[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
X_267_ net4 net3 net15 net16 net6 VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__o2111a_1
X_336_ _164_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__inv_2
X_405_ net20 FLSR_instance.flip_flop_instance\[28\].in _003_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[28\].out
+ sky130_fd_sc_hd__dfrtp_1
X_198_ _084_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[17\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_319_ FLSR_instance.muxes\[12\].input_a _156_ _158_ net11 VGND VGND VPWR VPWR _061_
+ sky130_fd_sc_hd__a22o_1
Xinput11 i_wb_data[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout19 net27 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_421_ net25 FLSR_instance.flip_flop_instance\[12\].in _019_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[12\].out
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 i_wb_data[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_23_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_352_ _165_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__inv_2
X_283_ _068_ _134_ _135_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_266_ net3 VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__inv_2
X_335_ _164_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__inv_2
X_197_ FLSR_instance.flip_flop_instance\[16\].out FLSR_instance.muxes\[17\].input_a
+ _078_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__mux2_1
X_404_ net20 FLSR_instance.flip_flop_instance\[29\].in _002_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[29\].out
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 i_wb_data[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_26_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_318_ FLSR_instance.muxes\[11\].input_a _156_ _158_ net10 VGND VGND VPWR VPWR _060_
+ sky130_fd_sc_hd__a22o_1
X_249_ FLSR_instance.muxes\[26\].input_a _115_ _111_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_282_ net5 _108_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__and2_1
X_351_ _165_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__inv_2
X_420_ net25 FLSR_instance.flip_flop_instance\[13\].in _018_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[13\].out
+ sky130_fd_sc_hd__dfrtp_1
X_334_ _164_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_403_ net20 FLSR_instance.flip_flop_instance\[30\].in _001_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[30\].out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_196_ _083_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[18\].in sky130_fd_sc_hd__clkbuf_1
X_265_ _126_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__clkbuf_1
X_317_ FLSR_instance.muxes\[10\].input_a _156_ _158_ net9 VGND VGND VPWR VPWR _059_
+ sky130_fd_sc_hd__a22o_1
Xinput13 i_wb_data[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_179_ _074_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[26\].in sky130_fd_sc_hd__clkbuf_1
X_248_ net9 _106_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_281_ _133_ _109_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__nor2_1
X_350_ _165_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_402_ net23 FLSR_instance.flip_flop_instance\[31\].in _000_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[31\].out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_195_ FLSR_instance.flip_flop_instance\[17\].out FLSR_instance.muxes\[18\].input_a
+ _078_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__mux2_1
X_264_ FLSR_instance.muxes\[31\].input_a _125_ _111_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__mux2_1
X_333_ _164_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_316_ FLSR_instance.muxes\[9\].input_a _156_ _158_ net8 VGND VGND VPWR VPWR _058_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_247_ _114_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 i_wb_data[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_178_ FLSR_instance.flip_flop_instance\[25\].out FLSR_instance.muxes\[26\].input_a
+ _068_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ net8 VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_401_ net25 _067_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[0\].reset
+ sky130_fd_sc_hd__dfxtp_2
X_332_ _164_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_194_ _082_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[19\].in sky130_fd_sc_hd__clkbuf_1
X_263_ net14 _106_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 i_wb_stb VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
X_315_ FLSR_instance.muxes\[8\].input_a _156_ _158_ net7 VGND VGND VPWR VPWR _057_
+ sky130_fd_sc_hd__a22o_1
X_246_ FLSR_instance.muxes\[25\].input_a _113_ _111_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__mux2_1
X_177_ _073_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[27\].in sky130_fd_sc_hd__clkbuf_1
X_229_ _100_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[2\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_17_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_400_ net24 _066_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfxtp_1
X_331_ FLSR_instance.flip_flop_instance\[0\].reset VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__buf_4
X_193_ FLSR_instance.flip_flop_instance\[18\].out FLSR_instance.muxes\[19\].input_a
+ _078_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__mux2_1
X_262_ _124_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_314_ _157_ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__buf_2
X_176_ FLSR_instance.flip_flop_instance\[26\].out FLSR_instance.muxes\[27\].input_a
+ _068_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__mux2_1
Xinput16 i_wb_we VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
X_245_ net8 _106_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_5_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_228_ FLSR_instance.flip_flop_instance\[1\].out FLSR_instance.muxes\[2\].input_a
+ FLSR_instance.load_seed VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_330_ _163_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__clkbuf_1
X_192_ _081_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[20\].in sky130_fd_sc_hd__clkbuf_1
X_261_ FLSR_instance.muxes\[30\].input_a _123_ _111_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_313_ net5 net4 net3 _128_ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__and4bb_1
X_175_ _072_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[28\].in sky130_fd_sc_hd__clkbuf_1
X_244_ _112_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__clkbuf_1
X_227_ _099_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[3\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_260_ net13 _106_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__and2_1
X_389_ net23 _055_ VGND VGND VPWR VPWR FLSR_instance.muxes\[6\].input_a sky130_fd_sc_hd__dfxtp_1
X_191_ FLSR_instance.flip_flop_instance\[19\].out FLSR_instance.muxes\[20\].input_a
+ _078_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_312_ _155_ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__buf_2
X_174_ FLSR_instance.flip_flop_instance\[27\].out FLSR_instance.muxes\[28\].input_a
+ _068_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__mux2_1
X_243_ FLSR_instance.muxes\[24\].input_a _107_ _111_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_226_ FLSR_instance.flip_flop_instance\[2\].out FLSR_instance.muxes\[3\].input_a
+ _089_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_209_ _090_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[12\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_190_ _080_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[21\].in sky130_fd_sc_hd__clkbuf_1
X_388_ net24 _054_ VGND VGND VPWR VPWR FLSR_instance.muxes\[5\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_173_ _071_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[29\].in sky130_fd_sc_hd__clkbuf_1
X_242_ net5 net4 _108_ _109_ _110_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__o2111a_4
X_311_ _130_ _128_ VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_225_ _098_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[4\].in sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_208_ FLSR_instance.flip_flop_instance\[11\].out FLSR_instance.muxes\[12\].input_a
+ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_387_ net25 _053_ VGND VGND VPWR VPWR FLSR_instance.muxes\[4\].input_a sky130_fd_sc_hd__dfxtp_1
X_310_ _154_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_241_ net5 net3 net4 VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__or3b_1
X_172_ FLSR_instance.flip_flop_instance\[28\].out FLSR_instance.muxes\[29\].input_a
+ _068_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_224_ FLSR_instance.flip_flop_instance\[3\].out FLSR_instance.muxes\[4\].input_a
+ _089_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_207_ FLSR_instance.load_seed VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_386_ net24 _052_ VGND VGND VPWR VPWR FLSR_instance.muxes\[3\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_171_ _070_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[30\].in sky130_fd_sc_hd__clkbuf_1
X_240_ net4 net3 net5 VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__or3b_2
XFILLER_0_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_369_ net19 _035_ VGND VGND VPWR VPWR FLSR_instance.muxes\[27\].input_a sky130_fd_sc_hd__dfxtp_1
X_223_ _097_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[5\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_206_ _088_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[13\].in sky130_fd_sc_hd__clkbuf_1
Xwb_lfsr_28 VGND VGND VPWR VPWR wb_lfsr_28/HI o_wb_stall sky130_fd_sc_hd__conb_1
XFILLER_0_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_385_ net24 _051_ VGND VGND VPWR VPWR FLSR_instance.muxes\[2\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ FLSR_instance.flip_flop_instance\[29\].out FLSR_instance.muxes\[30\].input_a
+ _068_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__mux2_1
X_299_ net11 _137_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_368_ net19 _034_ VGND VGND VPWR VPWR FLSR_instance.muxes\[26\].input_a sky130_fd_sc_hd__dfxtp_1
X_222_ FLSR_instance.flip_flop_instance\[4\].out FLSR_instance.muxes\[5\].input_a
+ _089_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_205_ FLSR_instance.flip_flop_instance\[12\].out FLSR_instance.muxes\[13\].input_a
+ _078_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_384_ net23 _050_ VGND VGND VPWR VPWR FLSR_instance.muxes\[1\].input_a sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_298_ _146_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__clkbuf_1
X_367_ net19 _033_ VGND VGND VPWR VPWR FLSR_instance.muxes\[25\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_221_ _096_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[6\].in sky130_fd_sc_hd__clkbuf_1
X_419_ net22 FLSR_instance.flip_flop_instance\[14\].in _017_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[14\].out
+ sky130_fd_sc_hd__dfrtp_1
X_204_ _087_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[14\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ net23 _049_ VGND VGND VPWR VPWR FLSR_instance.muxes\[0\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_297_ FLSR_instance.muxes\[3\].input_a _145_ _139_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_366_ net19 _032_ VGND VGND VPWR VPWR FLSR_instance.muxes\[24\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_220_ FLSR_instance.flip_flop_instance\[5\].out FLSR_instance.muxes\[6\].input_a
+ _089_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_349_ _165_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__inv_2
X_418_ net22 FLSR_instance.flip_flop_instance\[15\].in _016_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[15\].out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_203_ FLSR_instance.flip_flop_instance\[13\].out FLSR_instance.muxes\[14\].input_a
+ _078_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_382_ net23 _048_ VGND VGND VPWR VPWR FLSR_instance.load_seed sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_2_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_296_ net10 _137_ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__and2_1
X_365_ FLSR_instance.flip_flop_instance\[0\].reset VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_417_ net22 FLSR_instance.flip_flop_instance\[16\].in _015_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[16\].out
+ sky130_fd_sc_hd__dfrtp_1
X_348_ _165_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__inv_2
X_279_ FLSR_instance.muxes\[23\].input_a _129_ _132_ net14 VGND VGND VPWR VPWR _047_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_202_ _086_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[15\].in sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_381_ net22 _047_ VGND VGND VPWR VPWR FLSR_instance.muxes\[23\].input_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_433_ net23 FLSR_instance.flip_flop_instance\[0\].in _031_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[0\].out
+ sky130_fd_sc_hd__dfrtp_1
X_295_ _144_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__clkbuf_1
X_364_ FLSR_instance.flip_flop_instance\[0\].reset VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__inv_2
X_278_ FLSR_instance.muxes\[22\].input_a _129_ _132_ net13 VGND VGND VPWR VPWR _046_
+ sky130_fd_sc_hd__a22o_1
X_416_ net21 FLSR_instance.flip_flop_instance\[17\].in _014_ VGND VGND VPWR VPWR FLSR_instance.flip_flop_instance\[17\].out
+ sky130_fd_sc_hd__dfrtp_1
X_347_ _165_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_201_ FLSR_instance.flip_flop_instance\[14\].out FLSR_instance.muxes\[15\].input_a
+ _078_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_380_ net21 _046_ VGND VGND VPWR VPWR FLSR_instance.muxes\[22\].input_a sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

